PK   DU�Xx�*�  �     cirkitFile.json�][�۶�+��j�UҾ�9�@�M�>d%QY�^{�,'M���C�ZۺP�0	phc�3Ñ�q�㈒?���7�|[��]��&�!bܫ���ΏF��ڬ���}���{�|z�a�}x�n��Y)�҄f*LD&B.Eb>�<�2��4+�	n��-��Nq���q�N]��%N=Ʃ'8�ԨO)G�Hh��0��y\�0�	cEU!Ӽ$��3G�L"L��5�t�Q]SL��5st]Ri:.�P�,y�e��I�\�"����#/8r��%s긫c\��N0gMP]��J��T��
�X%!�"3Qa��$Ӊb�T&�c22Pl&E�R�̥�c.=
�9M)2�Rd.��	�t�IS$C��!Qϰ�z��0	]��.s�	P���ɞA)癛~�>k�5Ct���Ԋ����\ѵ�B$�k���'(H�=?A����d����_c� ����p����E"�k<L׮�
����Qc�Z%+	�=?�Q]���0#<��Z�pb�6�˱��o��Y~~�ڿi.�Bz�¼X�^�D^�/V�+�+�+��
�#��v�J��e���2DLa̴���EJQ޴��,��(ƌ�i@� � �y��L�aZ*�r��ĄEyӢX+�	*v�	5�S$�ʩ�XN(֚P�?(�~1��i�bs�1(���������'B���O,f~P�����(.2����Z��wZZ���*�|��|�i �v���^�������	��x�B.�Z���Т�<��O�0�2OӠU��E�B1OҠņy�@k�lZ>8��S%`רFc+�oj�FV�V�+܋�ȋ�Ŋ�b%�b%�b%�b��$�g?������4 ~L�@���0�b������H�����S?(�~PL����A1��b�����'B�����3?(f~P�.�\	�[�>p% o�"��� ����W�V.�\	�[��p% o�"^�� ���xWf��+x+G\	�[9�/����#`U7�.��U�w�ǵ�u��6�m]�:�y�}�"|Kfk;��c�F݋���n��:^����������] �����ӵ�0]KT�
�3jV;�0�J��1 o7�a�@���i��L6U�b*��3N~��zg{Gy�M�x���6��z�M2��"�|��ﾎ���y��P@|� �H�`�	�,?�{��)x�leփoBZ�`��4��$F�ž�7�o�28�&�Wv/�
�� �ϐ��!�R_"�c�~�Էw����#·�%�}{�$A�����"8v>,��m�3BQ�xl�dۍ{�g�R��TDF�tlL�ؠ�n!���C�0M�q��aK��7��S��X�2l�eX`2,0�DxE?%�p�+ �x{ ,ڃ�	��x����#��w`����0�3A�C �?��k�����m``������4��``α� �(�s�4�����
�ޠ�y#����T���;[,�Dr��)mx�1�"��h1b֎�������-!V�Xyb��&V�Xyb��h�h�ݢV�Z���j5�ՠV�Zj5��`V��.Yf5��`V������A�pcϰu|p��34� `�7d��F"љ��q�aV
2�T,4�Bvo����;���2':��Tq��$fHc�C��d�R���2����э�����(��^�����[��l�zC#r˘,�ޒ���2��ו"7��s#꽭���\�z�-r��8��^q�ܵ1�ĨW�6r�9�%�ȽcV�z++r�ǘT�^T��2�$�w�_c7_�U��6����_u��Š�tMd�D�&:nb]7񮉏�D�$�M�k�㦸k��MIה��Ү)5���AƗ�/GK5�z��j��l�j�ͦܮ�ծ�C.��DAe�bn菈K�M���4O��p��Vt�{��f^E��G�i���LD�������D�$,�H��d�Hf����Y�weC����ã�3j���j,���zSou�T��d���vW5�	��-i�$�t�`L,#���wG�1l���0צdi��8	#��E��B�PXH�(�k��#<�d]��7j����"�֕�����˫:_����4^���/�Sw��9�K��4bGK�X�Ґ.-{�t��;�c1ڷFb�M#�X, �R	��,)�b�!�"�ڋ&�11P�01q����qy2-�����!/�x����ۄ��&�&�6���ڄ��&�&�6!5�	�)�M�M�lBl
e�ҥ�Y�ܵQ�y��j{�Y�pn2��O�eB�4���d)� G���a�,�ӘFe(�T���$LM�E�kAY,�"��d�A%�a�_�~��Ib�+x@JJ�<1g6�̣x���k��v$:W�CNtf�c.s�s��@�ى'�����qc��cm$wM]mޛ��Q��m]�zo��$��j���̧������Kc4�)-W1�;]�Q�l���j��}Uk��Ɛ!��ٗ*o����z?;��c��z_5/^m���1g���?C$6"�ς��3+*f_�.qQ$	˓\� dxh��o�YPW����@$�R�@j��}���3;;.Ύ˳���q�J�"s���3C�$q��t^��~��۰��D?��p���Z�U�鬏�c/gG�n,/�EF��EP��ǗOC�������7Ǿ[%�M�������x���Ω�3C�ө�P��'|R�����Ou�$u�̚�+F���3�qf��r�i�V��I��Ɠ��5��3�^n�f��/~����Oq�Ah�
aV?�����ϒ�&Drθ����ͤ�<�f��iX�eZȵ����J�L M�MP�����G�7���eĿO����~�o��yK#ʨL�28�f!{(U�0+]j�3Z�$O�0%yAfk��\}����W�>�Id�'�(��gd��(a��N�S�P�f9�͟��?+��
�2�_����T�%iB�0�>N,����	M�QK��Jf ���g[D��h�e�}�-b)I�ޏn�[7A�.MXL,��Xͽ9$S���c�����S�L͂Ī����tn�޺W��.~:�/�Ժi>�Q��GmY��mоB�6��}z��m��5�B�f�m^m��o��������ۚ��Ƿ^}3��Ͻ�me�j�[[�ooo[0~]��o���Go������~Q�
,Z)v^� J>-e2��Rd(u��6�b0� �v<?W��e ]� ?׸w%�څ�i�����p��9PNc��"Hh�i`^��3���_d!�#K盯�B�[X�3D/@)"����WݠR��rxöW I ��$��� s@�R�D�R���UR@ ^��@���o 1� b> O�`���"<��-��WItxg�OnC�qrE��7_܆<+�����K�or��1��Hj�W�����+���y�Ƴ��5�R�t��Cc,5���"�����+"�^VD�4#�� J��8��H�Ai���	�����0���;$0��h�_� ����0f��T��]���1U��e�� 3�k�CBC@V1@���#�ih~��~q�и"h\�7h<+jH
 }!O�T�������aA��{\wP�y���;:����-Y13���41����~���{L 4�<�~@�j����CN���&����?�����b�^�.Q��+��7Q��K��.~Q��Z��}x���m�g��PK   DU�XK���(  �(  /   images/1042b8f9-2e87-4dd7-a644-1e53cbd80f37.png�(׉PNG

   IHDR   d   R   ��q�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  (|IDATx��]xUղ��O		B!Bh����ł���P)*�x�*łPEi
�"* E� ]Z����s����t��y�����ee���^{��Zk��ʆ>|�/�|x���ʀ��>.󱛏5ο%Bi���+|�'����Z����A6��Gh0������A�V���7i4Unn�'��4�1|l�c�n��$��tvVԧ�~�@���ΟUd��)22�֭[K?��s�ڳgOz��������D�o��o���J��N�#������o��իW����n%����5��o$�R>�Acʔ)��c�Ӂh��/)=5��v3� :�5mM3f�,�^|�E:v�X���]�6���kԦM!�ƍ�ڵkG���'�VO?��m�aY��TvR�t��[�z�H۶m�U�>���~��U>�xV��+Af���h��kגV��_C�5�*<��;�`�S3Q�Ս�b���'R��.�a�74}�4��uez֬YԼysQW��z�A o��&-\�E�;H�#�i@�F���Lb5oc5�M�o��֭��&L�N=z��aÆQ~~> ��)$HOr��#11�֮^L��مj�� ��ʄ��[,�4�C�&!��,�!?Eƍ���?���lڲeK���ر#�����W��IKK���p�]w��sߠ	�GSXc#�K�8��,!f�JU�ǧ��oﶔ��C�M�a#����>�f9��^� 0઩S��d���#?���l�wو�d2[����%%�ύᇎhь��U�6�Ez�ͷ`���'�,4������#΀V�a�}K777���+��_H��	f��.\���Xp�,ԭ[��{o��{��> &���o������s��c�����;��$wwc#�v�x��8뭷โA�~|�G}���h� KĞ�y�ѠK��U�P5�/�d0h����XV��6��\;B;vlg��8 aaa,Yf�O�>}(66V�j��;���x���{��ǇN�:E���>m�49g2���W_���S�~�(==��S��s���O?Mk֬)t
Ч��B�o���Ξ=K��>�5J�)�#����˳�����6l��;w�4A0�_��<ځ�������A����_j�j1�[g���3{ǋ�A�~D��9���Z� ��<#F��� �PS,W�LC�:mn���G�^^I��=��A�����L� &��ݺ���?o�����;�̃�*��K�.I\�����p�R#*���������w�A-[��ƍ�'�|B���;͜9S�شiS�"�^��Gy��}�Y���Ç�`d�8l޼���
���<�w�3� 7P����S�Ӡ�[� �7]�U������2��w��{s��Z^��ui��Q�����?�����#?�ԟo�~�j1�V�}��Q� D�%����W�@�x�a��5�`����~�^O���y�Y�&���#�p��U��'
"�����Ӑ!CD��B�xp3���+���ôu�V����F�Qxx8}��wԭ[�BUI�.��\�B�1yxx���ۅ(�
�S rrr�p ~U c���#Ow+3�*sTZz�O#i��ƿ�aa����^�1����1J`�6�q� �޽k;*A�> H#p��G����&����]�����Bb��S?���fb���ͷ�C��󡨨H1�x �̣�>J�z���>���]�&./�P/x.��8r�xi���؁1cƈ����rr2͞=[	�P�V�Zt��!J׮]ŭQ������>0 � l �Y��u�6������c[]Ｚ�>t��׊��9w5�{u$�N�m��L���ky��S�
�v3q����f�0�l�$k��<��Ru��%���%p�?,#=��ԩ#�:t��z�)��E�	�Ce4l�P�>�]n�w�.���p��m�&�R Tu�X���p���B��n��"�W|�|�]��Ni�����+�^\.z{4�ך��k3����q܃Lw�L%/�+���LA��%dƤa4�ݵ%>���É��9V��{ԪU+AR�-DE=z�֯_/z��733S��ڵKw���i߾}b0A����"�]�dI�AG�	&�Z���9s�3��� ���d�IK�.��PY.��w(�/ #�k��Ы�.|jy�z�/p�����^� '��ŠVB��^�)�����"�3���"Y�1�1��ʥ��z����* 95�"�s���BCCE�aG��@"��U�hݺ� _H��4�;w�سO�8Q�������/����ʒ�` �k@��dʃ���{��"O�J-�ݙݽ�A/]N�LuU�k����ڦR����y�&�9p�� @J�>}��[��+WORx��Љϱl�OL�E��Ѕ�Xz�f���W���LL���j���6�K̦�a�iƾi4h� CT$a?�y�@�#@���F��>n�xZ�*�����I���0#�[s���s>���?s/��@UQ�Z����,���	Ԃq�_�Be���_ӼwޥY�~�L��=�5L��t[�ϔ���;�|}<A!�z~�-��4�K�c�a�6̭It��e����h�N@�^�Zm`` M�4�Pe(�@�� ��	U�$��I�r�����R��X'55E����8j܀}|�r����.�h��W+&A{PRJ���F�)K�=x�c�ЫoΠ�/M*�o!Av��M�I�R��J�I=���+��%���[��K����-�m��_�/�eb,ᛷ����E}F�'�$�[�l������v�o�0�@����_�>M�>]� ���ԩ��Hl�b?@(�ָ?�EP��O?���ɓ'��ŋ+L�� �ȼy���	OP`8Dm'�1�Ƶo�dW�X&����e�#��r*���L0�w��8���/�m�iS�ґc�C��H�T��̖�d�h��3�vd���o�n�7��/� ��4@����+����@��/!;q�$� �( 8�T� "zxx�<==�9 "�4~CP	�VU����ǎ�N+�ͥ����Z���<��q���0�0����eܦdyҤO�3r{�{!��رc裏>�@��~�~�ݽ��zv�Q���Q�Ё×���3%27n\�_�)=�P�sp]�UA�A�����2G&A� 
���zO ,�)�;w�iH<+�B�ѧ� ����,�`�\��1�B��V��n��1�'|��,ں�y�5���ͦѣG1�/�_1�1����h��RTd�[�9YM���ϓ�Rbփ9��a��-;��K^��D�h@~��`��r��@E�5i�D�M��p�
�|�A�xxw�O�i�z��	�@h�--�YY c"�B�`ђ�i�ʏ�͇��[G�}<�0jQ�)٤��Ґ�'���Lp��M*Pb����z��O�2�Ll#._���HN��� �t�"=��Xڻwo��\axb;v��EI� �D��)V�ZE������8�͚5� Q�@,�<D�#G��{+��� 0"�=rg`�G}�	��k���ܸ1�3}�j�ɑO�f�B� ����' 	#�t^�ϯsl�$���Õ�N@�/�g�3C��_Ib���p�xs�"�Pg�"(N </���A�3CZT� ��O��X<���dqmO�<Y.#d����H�"����?�˒ ��� ��q( �T��;�P�
@E�&�p�q���z��*A:���mى�3,�>��������Is���
 �ڀΝ����EX ��'Ӝ-��m�8-�Q$�K��[q;*:^f�Z�х�� �V�]�At�r"{/E�檛7���� P����l,7m#��O��{N����8PS�IVYGODWۀ�ס�/?O/�X �	�)3��͡Yܞ>kۆnO���,��4i�zu)�'$��h��et-6�f����Gt�j͚>��zo%�q�"σ�u�O���NƺY�ڇ�k�"�b|�a:%F=��5�L�N�!��1�`��bұ����O6����5��,�`�Z�q�#n��D�5R`���7|�\k�6P�OH�c� ����J�KA!�Ǹ��,
��/��&m��+Fn���Ƶ,�	��NF��+W`G@�B���ͽܾE�����b:��G���ׯn��u�ۗӔ�k�8�icj�6�BZFPj���L��B�l�X�>�&��qO��؅��Jۮ�q.2�٭Ζ�>α��v*)�VI0�*A��1`<Vk�فrgj��{�r�F|����~tl�~
�W�4ZGpeb]m/0R�>R��]uj'�B#�f��f�aE�ʥ���Tw*U	�o�VEER F��}"Ƞ�F�)�bbdf�Q�.aԥC(<r�Ծ��.\�8�2�,)��2w�Z�9ر��l6�ߏ�N�1q
��b�s�
d��h�6���}�p>�T�?���_�<����
�j4�龻�QRJ��߯��
��J��/��A�V&`�����#��E�d��~˖-�Z��E�.嶗W-،�!��ߛ4i*}��=(4�-_��D����C	��jIGD��*#Y	>@j��5�
�51"0��Zvz�z	r���C���d58�� �`�FJ����۵��<R�J[�m䤐�G���O?�DC�Jz�H����o��t�x
m��2��K � K[�n��N#%+����t�¾O�9G�� ъ�wM!�L�炴�rO��(�c,6C�%��4wJJ-��Ĳ�`�%tu|b:��<J�i-#Ճ̆:x�ef[Ġ�5�Kލ|i�敔�G�9Y��r]C[� ܷ&��r	r��:z�<5k&`�5��:_
m�]�, w7:~>��|���t�_ ��Ӡ�(�邖�Һ�h��=ɨM�Q�����D��e���_v��Ke��߿�v��N"؋ ���͛����W���`6�G��eɲU�0�*V߹���Nm�4�<A�����&n��{��1.i���Ȣ��"��Z������	�:��l�;�����?��p}�f���eA����E�G�#y�:�B9B��lZ��6���S�
@j�{nu��^8�J�a6�v���!����,���Z5z�xY�9��"���m@�'Ӻ�eo,� �_5j�O��#�PX����'��_~�ܗS�0[�jޖn��_���H{m��V����+q7�¼� ?��lv]1��'��V��3Kp'�\���}�� *:|2���E���rK�Z������N��+.qzZK��.]I�:���^m�\��]�f�%KD?�j{��Zu�%
o¢�˶=��y��M�BQ ���`����6��e���
�Vk(%9��әT枴nS�kJ$������n#A���Iz�Y�N���gCm+�8&`<iƌ�@��ŋ�O �y� �dk[͠�s�K>��6Pp�ze�-� ��Fz`Pw�!a�o���L�$3v�l�Q�J�ϮQ�?p���̕t5�˂�h�~X���̾%	�Դ,�!�/]��N�]:�̗
MW(�.������ykd�
V�#�R(���u���?�諯)�o�1����\6�P�i*�$)���RR��+q���E!�qw&�pd�8�� �;R`.!a)���<�@:��8�Pu}CO��F��&O�^Vԯ-��Ҳ��^G�	��(8��l�/V
�T��e9ԧ�t��B���E/O*�aÐ�ܚ]�4�=�M���,�n��<3v؏rs2�Ա��a����w:w!�0��䟀,eZ�:���F�&&�:�%+k����&%���{�x+����R��H��Y��_k��Q@@��7Q����T/o_
jB��t��4�:%=�D:��1Ee!��/Y<���~]�l5Ġ0N��pג��W�}K�CV}�C�nI����JZ��j	0�>_A���B��� G��<C�~2 ����GU3�7.��GǑ�Wm��/K�7PZ���^K.�oɑ:G�{��*rө�;w*Q̀ ��۷��\qXX�Ϊ{�` Ż��ɧw}KS�N�\VM񲰚���$����̾���ի�c������z*�����?i��C$*{ȱF������t�ԙ�+�N�(��=�N��v��O�>�nmu��Y�`�{۶m�XX�
���5qBE4B��.�	�r����ceَC����h�hQ��B�ۄPߞ�����^VAZ�&Z��}z������B.���|������iԨ�+�ǎKW�^��|z����bt4-X0�Ə� E	���a"�=s�>�`1��Ҕb;u�lŋ�	�/&��?~\�IiP!����5 �ޓ":���Gi��?R������ɦ�����
nN�}O6K��D\h6H8���b�D%+"akmi��RΫm9�l�wM�y��G8T����d�?���u����X�r��+msS����dbψ���݀}�Ӕ��Gu|��n�^�������<j�燩���9A�\��X�e�~Hy$���"�����vE�����yw>����\�aw]]�!�Z��l@��JG�y�c�t��e�����{���>�b�	2d�T�=z�\[�z�J-�@l�%��xq-������/V����tѶ��ߒ��v�����l%�=Fw�3))9���$-Y��Z���ɦ�<�tAF6���l���(�E�o,��h��1;q�z�(���}��6���j1	!���J�ö�T�+=���Ӫ���хr
�Myt����C>��Ξ���I�^ڹ���9i�6�9�*�_8���"���ɭ�N&����̢e7�￻�I��kD{������o����O�=]�����R��ftp�Wd�ϔ-��+5HEy�����:�E��Bi��)R}бS�7�mJJ8O��l����+1�U6���"�#C,�"G�U�p|��.�]�M�i��Pbr����Iܶr{*����$k;u����%\9Mi�ژ6�JI͒��鳗���"`w�v�iU|�C��P�M3SJR���k���R��ܹ��
dG ;1v-Y����u~~~r���Jm.w�biP!�@��ň��b��@����H��UŚ-�Z�,�V�]�����꜋���Ħޯ������Jn���ca�����bYڴ���ma�����{b��Ƒ�Sd0!Ω����<��!ԡmJHʠ}�)���
d�޿�ԙ���k6lC
��\�O-�nzvmAV.�5��n�my����2ғ����,Q�(OŶ�O_ھ�JJ��\V��a��q�X˖�J���bcα��ei�),t���D�.�����}m�����@z������y��k�//�Av�����rr�{�n?L5rr
�]���Y��a_$�2,6-śԴc�^����;9]-^dYI΃G"���k��昖��ʧ�m���gNҁ�D]��R���S�:wh&���_�����?�,�o1�'��MH*Y2������ϫ�J���9n�#G�3!�FT�S�r0V�d���~IjAJ+�W�R|e��@y�������`��'ٍ��6�SF|}�ng�l6�c�=/� %�rQ��P�U��0�lEq�9�V�ݻ�Th@�E�po�*S-�F��B�T1�~C�gGmL����o�7C�C�ŪZ��rT �K�.�.ٴiS��4����ϲ+R���V�\����R�܄ �w�T����!����Fӻx)U�ր��fp(�? )�$��x
U�p/T?Ey@���T��H����|����hIP.AU�����i���P2����駟RU �bw���G�Hp/vF���ʨL|!��rM���k�]�pA���yX=��Zպ'�G��ؐ��[���}\��U*dCP��-��m۷s�m�k�b(..��
  �t:�&Z,6ڹs�����-,��Խ� �����N0=�(;(�������!Ծ}��@UmJ{@J0^ԏDU�#G���=S�{U� � e�{~N��t
��b�MF]K�{�L��m��Q���Y0�u���R��P�Z%�{���m;˂�+גh���왔�����MJ���D�k�}�qYt��n7BA~�A�G�!������ҙ�U�FR/k��Bw�d�E���_~�Ev؎|�K���⳩a�]�I��@����MK5ُ��l)��ku��kD+V�Z�(���U�J�X���nڠ��u���-f��蘑wP׎aH;�rZ���ݽ-�dK�z���~��(��?6zJ	��-yulJ�~'�Whވ�}�.!"�=�C	����ۆ҇�n-�� n����шWfOV�Uu:�oF�~<@�m��H_ج��U���ff4dF�j�׻G�賟�艢E�ʂ
/2bh_l��������&�����^�[u?u��컮/�5m@��삨�R���$������������9w��@�vj��d�HH�����F��8׽C��%+�sr>���ɧ��n:����e+��^�vi?�{�9 �Ȟ�{]�^���9 �B,���ha��<F".//�I~�Z��=�%�S��<v\�@��-�<���E���b8Ƹ����q�v>:V��Z	���[����i�F���u�?;�չ�2��3�&k5��sڭ�왞n+ڵiR� �X�Ks8���j�Ie'7���߱~��#�6�_(%(Q޼!\�ϼ�t��ycD4����q���TQ��pD˸��9�/܌���ԨU)����`������0y�c�ɒ�ձT��l��c_�ws%H'�J��f.4Z�	A��V�L�6������Jߛ~#Ad����(��̙E:��.b�G��n�b��-����H]Xm���\w�&�� ��蟞�o�'#�i$)ɗF������@�Ǭ��E���� ���+`��F�����]�.��&�U�"��r���=���1(Z��`c�Z�z�ծ��������g�2��T����������!�(�'j��bQ����=pO7+$���4���{C�5�Z�s��aO�\6�޵<PDx�1.�a��q	iPA����A��0����0�0�����_�I������=--��ݷuwmOO��IxNa\�{p\0�jL҂�@�|�Fk5���x�k�c���,����B2��x������Ú�����W��o�ဆ��0��� � �qoY^O�w:��E$���v���/��fx�W8p��V�fb4`n���P���c��cQE�o�yL��1�~¢ޕ9�Jà:������y�u=�]<����k���27~����H���0� �E��>=Zu�{�䱯�[���Y�1w�g��v�vTw�ُ��[n^~77�C(e��P����KҐq���֎��8z����w�� �� A �~��L*�+ۇ���:�������w�Yy�t�9b 7�������ᚮ\�Mvi�t2R
���`�;ѱi��n�i��%=� �Ut���X%��!r�
h�փ��=�JX�wu7�B���f��o�� �m��ȭ�4��`�Z7���S{VVQ}�j�xj�k`�}��x�p$}��+�A|yr9? Y E����Xf@}_���_���%�����ԬI ���eAx��f��Mg#c(��æ`�����-~��'$��s�ЁAJ,��賭�nץ� _��[��5����-�q���D]�+�{R ��T(�ǆ'���K�
���� �N>���P���9*x�� �2��@�҈P��e��8`��
�/!p� �;�w6�^���A���8�g�bK#� d:Q�ky�)!��D*�@��oUrG�P2��/�T}����H�`j��ue���2��"�T)�����B*�HV"{�t}uavp/Qqa��g@o���H}�/��@"�	��G�ߪ|� ���1��G6����J�A0�_�8 0J���Y�2�HT�z62��L�e��=�#���������&@�W�W�Mx)�7#��tU�{"͍I  �E��$�}*�0 �w+�3G`7�__@�F��j�`��C�|��:9>Z����;@Ea U�@LaFdq�<�� �:0��)�+pP��2ҘL�کL�&\UI �`5�1���R����|A�jj��?���B����M�OV���a��&�T/ s�J}un� B]����
7Jf+� ������V�&���x�@�dR    IEND�B`�PK   DU�X�;�i �N /   images/10c49116-c115-49dc-9efe-e8b38f603c33.png��y<�_�?��J��DQ�J�TH�%����$�2�s��4(d*2���L��<3;f���9^������O��~�庮��Z{��z>��neE��{���`0�eoJ�b0���GjJ��|�7���5Yuj��B}�{��MMk���wG�#u5��Q��wm����Xc���/<23�62�0�`neN?����J_Uw���1��躵6�����d�}N�}u�U�a���?VT\⿣`h����o��|O
m����c
���L���^?qlǉ�D�Õ���$���r{]Ub"���H]+�K��v}}�-�f�I������F]Y�n�/r*�r�2�=6��]�Yo�yy� �x_�V��F	�ln��̑��}��1s�g1��
:U��H�}�Kx1�T�3"R�����)�1���2V�_|�XP���8y�����{�����^����DY,�c*�}s%Rr}��uf�@o�r�{������6�i���9�KMmWU�p�y���92��1����%jA�%)�{��|��Ķ������vUB=�튙�?������i��6��}v#+���	�/�;�W*��s�4��I���ؤY<w9Dz�Ӳ4q/'N���0?hL�3��#g��
����u��f�z�3pL� � ?\�/O�4(�_6������$�zS�&��ّ�4�qIi�E.\/��9^#xH��x	<<�a�~�d�+����x�oX�����l�E�Ԅ��OP�=�N��)+Z�!By:�$T�5�;HAl:M�v��G.�_�#�>n�g�Cx� r�F`ҫϝmOj�M8���'U�I_R�'��I�˰[䁮���x�\L��4ڇ !�Z9~Jl?t�뱾eѰ�����{+'I�a
�l��a%ɣ�+)�xG��}�EK��{�"u#��������u�@vSy2������/�|�S��Baz��(I[4D���j��(�jm��m�:Q�"G'M��C�$���Շp�>s��$o�Q:|A4��/��&W,�u�F�f�q��l�q8`�7��H����t�=}Y�2�����D��8����m,�IAܞS�#��M�.y\�di�I:<1r�]��"j
��w#�l�d������Ê#zW��4����!��/%��	�Cp�j�'�=�i"�nZ����b�����W?��*���.OZi��ȱbf
"��<�����''�����6%(���O�7�Ԅ�S���l�С&�o/�[��S
�y����pj����O�6n��!�M,->�#e�H��;�|�ʞl�'�Y�|���=̗��A�E���b��1�Ge:�)~ި�N�����9g��k���˦��1�=��z3�d�s��g������չ��މA�Tj��F��+IQ�p9�=����r3�	#G�{ؤl�X�T�{�g�C���Z�4ъ�?�����N�77�i�9�i)1#q_b��(��^��������'��o�Ze�Ƣ��M�y&���g�j�����Ԙ�g,���@Uv6b�\�I��MБ&����b-������8%��vf��Z�?�O�$OWJU�cӠf}�<��W��c��3���&�S�o��D+��}ghi�#���	JLKJNNNLN�� �I.�B.i�ML�F��ߐ�������	���z�p�0a��{��u��BY���1f�X�7�����]���J


Ih��F�:�MM��s̓�u�V�}�2�
Hw�X��n ��������N�#�5m�#�_MLN�|}��f����7i�^<u@|�
?Z������F�k�&�N�������W�"Ѯ�.U�X�S>�3ϑ}�\ז�p�T}�b;�!���VBx�g�7
���ѿ��Y�uC�u��A|^�Io���[Z��;E�W��_b�Δ�YUU��Ř�'q���.���z�r�^�^=6VV�$.��MҢ�I�[V0	�i�8�}N�Br}��-�f��.�������!�?�~��7!�O�0�)P��X����φ�̏by813S ��oX�������Ʈ��N�VBdmb�(�K�tU��a�
�W�? �>Kt�-jDG����b�ڬ���	d���N����1�|]Ԓk�z鑪�0�OUUU�5���l'�*�jf.Mu�U�X�L0 �E���
O}/�jV� �]D������6?�4ޜP��j�	������# S�?)sW�,�'Z��+���p��ҟtf��X?�XhN}��s����d\���ۇQ<�#E/S�0�v"U���J�Ö����J?5���l=~�$�̸�Z.4�T��F��: �%�ѽ醕�����0�(Y���c��*0��,-�EF+�|�RS"��k�u��J6�VFB`����D��hq�wP`abԶ���*&�Ȁ��NMM2��;M~Kڝ�b}3���(�Z*,ZKLI�h(^��t��j��x/7gWK���y�$!���c0�pcgg�ӑG��f���O���DY����S�w�AR�رc�$=��~\nMs;\«���Y�%�:�@0P�%�ZQɨǢ�����O�v��˗.U׼��t���l��>!{�<:ʦ��_2���ge�w��g����*_��ڶ���`��o\|��͵pu"��(��LO�|�T��������iph�ˢ6���!�]���>TN��D9��J+N �V�_l����� �gTl�NHwc~�Q��T��k.��;���lc�!b���=}���th}�!�e�ۼ���1�#s�5*�:X����m\��������P��T���%��%�A���8v��ډ�s�����w亳�3Dg����X����od؎�m��#onbw��.6��o	pC�y�Q~�r�DI����+��B7�Ь��2�/�5)�N�+�ڴ\��&A�H�{��HZ�4#)��-���#!zl��V�f؎���������͵�89��b��=}<�Z��S�vy���%�E��]�n�3ѡK�v�u�X�V9� ��#�P�t9�d%�I��b���������'��V����a���ڸ;����0���創��MJ u8���B��cw,����}�^��>�/��B�W[�n@�o�Ἰ�h������i9��}@�4Q���6��,���N�q*jj����I���hend;���D!c����x���S�&#�I-�9�۷ � ���À'j9"��*�;J��$��f犰��m�x�\No����s�=�W,��pQ��f��$��[��j�Sj�Tܠ���k)U�������֗q�o�b�k��H�H_k�H-��^��k�,��_���&��N��|*.�(�\L�.}�KM�s��aB�����P�m�h-����`�����zyB�䘭��v�;M?��I�]��9�+�1������i��](ZP�V=��J�~�:�6tm���L�'���(����zye�u?U��?]��v�X���5o �tYH�Z�+2؉�:(�P�w�׭��'���Ь�ZgC��7j���؋��^^��v�$���Օ��~�N_����&�1i���L�`��[�	J�(������:_F��Gc���,ҐP�)�Q�H�;G����X����Wk џ�rM��ñ7na_�����EY� ��Dv���>8�����ڢ�A���hJR��oѥ��	r�1W����!y�L��R/ڵi�T�A�î9��m�i�'.$�ԫ���(��߽.��x���M�"P���j-�`,>���J^0�s�F��e��h\T��A|ݟj��t&�'w�a,��(�h�T�s�f	���IF�����ɗ=u�����6*�m>Iɵ����n�.�5+���O=�uo�bc�a�U'�|�j�?~Tm��ad����vdN&C�(�ͽ���a`˹��T��dϔ��s)��;�Hc��_��5�K�AK��c� ��X"�E�c?Ux$X-%�	����?���Mu�,�Z�I�:e���)`d�>�v�����L����y�?��:(:��"����y�dg�I�U���,WK�Y��rw!?�Hy�t�?����A��:��KBB	�O����a�a�Ϩ�KO�mG��]��W%)��A\�N��������	�yYޫFU�>�vQœ�;u����ǐz�tx�?@�Z�I�}���Z�ŏ=I&3����'O��PZQ|�"15U�B�����t��[7�������<�X��װX��;я��WN�B^Ӻ�I5vt�nE����@�[���׽�]�؞�%	�=W|T��!��4�A>��9��M��!�>L��/��MP��7�L�]N���~�:.�۷󢢢���~�ށ���$��$Ӷ����5���z��]x"���u�2��ctt���K7mOڜ����nik�����)h�P�o�<��!*��4q氒�۷o��?���:�P2o�O�}K����#V1;i99������4===�"�E���(��55���v^�~�%�a<3l��,d�2��Y���y��9ۇ0�����l�7���L���O>t�k��j �z~����(T���,�G�>|�4�5E�:�v��{]]��w�tYϟ?��D��3��L7��'�O�khȀU$�#:�Ix��CP@�iz����}AVœV8W��r��eӶ��
'{���ӊ@V1C3�+}� �
G&��8 �}@��ì��`�azA���4��df6Qy
��6|��h���h��P��d���ƣ��*����I�b/�OGBH�	90FFF���U�����׻�'��Nml��ʽ���8�H���eP��T���>��ﾹ�"p�#�js�}�y�"�-e��էҏ�:ø�.�G�� �PҲ� ����ؿwl�^�@�0�;�:�3A��ܱ]#���R^U^�GPQ"������W���n�i�(k�g�=�nB�4��ZZZ�r�9�����BM��mHx$�P�f�{����������r �2;X���1�#�քlt��A)�Ue$	����o���>�!'���լ��ӗaG��幐�'��_���.���t 5��\4K#̌�D���!� i%�'��YI����f��4����Qp�] I�t��o��J���Dk���9��!aP�Ќ+ �+~x�3�\_I���t���2.qԎҠ����{<c�3U�l�Ch~"���6&4H�q���4n/��,�7��'��_W(���W� W�y_���,3���&Y�GM_:  $���*|��Q�W�Ʀ��N�5g���O�yg����H�C��:Zn,�'D��SYP.���S��ىj7���A2l����	"�6�5��C�CAAH�@0"�4�r!+;���q��m�㍋R�[]�W���A/�Z��
$�7	ӛ�~!;�1�/���]��Å��	'�YD.�CՀ��0	n~�uv���z�}�Y)�d[���{�ᐉ��ڳ�V��֑�Hm��aY����	1��٠����h���@eig��+�����#9 8!�ڡYk��Y(�J�^,��b��%�5�ADx�U ΛL-��2W���?�(D�͑ŶE%��5=��_�t��&��|AN.�	���j��ڠe�6վ������Ǹz��)�hW;��F%��(B�d*n�P�֐x�s�F]ɺ��t��"͡n��<]��4565%���olia@r�^Q�L��ͻ���:��J��Dl��QUu�D�ʰ�f�ԋA�w[m���RyCA�@�u}LFr���n����ߤ>bll�&֫���O�~%���� >�M�-AV ���
�ĭ䒘��怔�|�qpk�v�Ӎ��֏�|�溯�Bd���_�)����ajj:!2�)u@��ƸB/�8K�ﺺ���Ө�vV�*�>!��dAl�6ޥ��̨{�ц�z�/QW��x���hj���@+牏���
�rF�t�jP�;DVokhh�
���*T���d{�߾�Å�=�%KrXD �)Ч�N�����RC����峋43�$�;܎{�����"��}�C?9�P��a��_�w%�i���U崒,�dҨ2���\oul��1蘾@i��e=?��	*�ӍJ:���KzEox�	MNM��}������f:"6/�
�͸/���,���+vUS�rV�4�r(@�
:,� �TW6O��D	�aqS4�Z����I*�7ڂ�1��.hX�ߴ�.�-u��٧�w�` I��Te�Y� Y#��C@S���.$�%���v>�b@�l�s��.�!m���|�+�8rA;�Sq�Jv��L������ڛ��E�a4<~뿿��u���[P��H ��e��܊�K{�{{���\��i����x+��@�����~>����:�.z��XNퟔ��c$�`1%ʒ�̎=/����.@lPU�N�aK�J�H~+�[&�ۨU-2�ʷ5���Th���v������K�� �����y��z[]~��%��ܶ6�ՀB̌z.�4L|�Ѿ�_6vvU���2���� �w?#y7X�7Ļ5��-�����~Ņ�N��1<���{��"}�w�ڐ(`�y�y�z�> >>�R���W�h�j�I3�b�o�[�$j�hPw��t,�2� �jY싓w��g�$�uN,2X}���r�� �AU�\.��,vqԶm�=;��u-0{��Su��<�=����&��KKKP4�<�V?������V*�0�����<����!��F�04�$�w��Iշ��	����D,Q�[rz��-�Ь��@�y 
���Q������Z�>�-D�inϑ�����,Kh�����[��h�o,΂�Ͽ�
�Z����W�ٰ�h������ጀ���H%Dj��y�A����:MԔ:9�����F�U Kˢ� ���Gv+ԝm����\��v<P�I��ƣò���р��т2v!��������ԛ���%��t'��j~������/QZ`��(b,�����3?++bF	��R�6
#\�:	M0_o+�C(�I���W�����g�\8%V�[��wF�;K��^w��d�\�}ҝs~1��%M�����軱�m�^���g���O))<��5�.��y{�r�܇s> ��~mm�����BM��=|��;��/o���^��Ms-jJ��n�~�%,���Ub����,��l�e��^ �`��p}�c
�s��<z+���Yd���bs~�����
S%%(�?��8��Aа�n�w��ϲ$#����pb��VkV-P̈m�,��B������t�����&0!Io�E���0Dt^3�2��Xk������a�	b�q^l�@'-=Y����n�K]��+#!Ϊ��{��t^E����Gx�����m���Y��e@�l^}AY	7#�j�m�V�/~kNPB���Nb���:��Dk]�i�!�O��݂b� BX`�j��7���HՌZ�wf
��}�����Jjz�)@ʡ�5��P@��T��wj�7�����ƴ�$�h~��Ba�W���z�h��jC�)���/~D"]��B�����IwY�[�ug�[�Zo����*H�x.6��)(�NUbh�KQrc�I�B���>B���.��}~��k�1b����Y�i go��ؐ�B
��qnI5��a�y��O�5w��R�Ӌv:0����s�g/�Z�'�|�W",���2���D$�...�(�g>�U�D���>�"��y�����΢]k$y; L�6'������o	��6�׍���w��Du%��7�7����˗/7��,!�N��:6M��z�m'�SR}?|��6�<̬��
WbO�S��$��h������惙�?:w��䐫�?��V���v~w[�Zx�|�/{���b���)C4k{c:o�B�Bi�\��/7��Z�2 QJy�Q�K�*��m�x�_�<�BO�VCvk}޲Ƕ�::�8��Q����I\9:W[_����oQ�����X�Zd,a"5���D�;��G�u��)�@�G��,o�C���2t�����5*��YލK���5o��,�/D�/2J�r^q�t��1�6�����]q5�R�hC��	����[(�Pe�����v����F��⎜T���0��(�e���ϟ��_�G�=B�bq%¾�1)�5a��DI �C��r�� +�5�b�7����s[%N��Fe(��W����J������ľ�RDѡ�D���Ԅ>`�?����o����f�N�!��NVNNU��+�.���X@��*�أl�	H"��'ZSԔ�{��/	
V�6�P�`��Z.��Gt�_jmk���q�+�F�5=~~(�d�)� 58�g����͝�G%�:й����˗+O�h�J�h�E�"�"q�t}ZD�R��~$��3ӏ��f���.aM��AAV9�V"�(7)>�-c����X�#W:yXh���&k?u�ˎ�DzA}�c:J�R!C�0X�SRb��D.���w
�%� ���PƉ3�>��)���|צK$�_ɾ�L��OLI��72w�|얕�U������\	M��At��K���$w!�� +�%j�����UԆr��;q�F���Ǐ��n�we��b6��Y�j��v�E��d���c��u�H�Ň��B[��<w�zk�]^���3��m�i��0�ߢ֫�Yٻ��9!����tB�hT���P���t�mmG�u�u��֧��Z7`s���t44�Lf8MCz�M�Γ���H��NϘ�LQS�^F�#MҤ�?�/�� ����q���[�� �l}* e��_��72�"%����������6���B�L@0�#���K�~��م�G)!n��$���J-�AsФ����6tjVzʰ����F����-��=���Q��Ȣ�������a��+!*C���ޕgm�^����Da�ɭy�w��[O��3*�F��0��Y(��{���I@�G�s�-��>�J��xS(�э���ϔE�����[HA��w��岔}����.��b\]7�%P#>sK�h_�?6�P'���_N7��B�5J8%��ߡ�`ۇ���t&��ML>�O����`��4�;&�nn���Yo��GM_�����\.�č��2"V��$bq��ɅS{#h�g\2y�ـ63ȿ������:�F{�W�;�2��+,�DZA��DKi��r�����ҝ'��fy���iV���蘒�P��w%�L�;�t�pA��k�������X�h|+dr�	�����5�<�СA*bw�GB �V<��qjޚK>�KXt���(sȗ��q
��p��JlW��a�]�#콩�-)��0���G�^�*�V;�.^���zOڶ/�Bǃd�ܿ� b.�u��(��G�s�B�as[h����������va�;= VS����t_I�&�C2p�5K	��R�E��#� 8�%�]Ξ?:�&��9O�A80m�;�l`�[������@��d�m|�z��`�H�}A��O˞���|	eiK���۷G��M]]��JO=,eѠ븩�ϼ��d㟹���߯���e/�L��⪋.! !�`X��8P��=�n!6�Z�^���b���uz���aޢՉ��C@�����-��C�Y�r�E��~HWucҦ�c��fؓo[S�����TEC#�����D��[�F�@�Q+���(`�|�/f%�9��B��ȴ�O�s*����S�@�I	������+�)x�~}d���w�+��䶵և0E@,*�^rk=��y��c����L���e�����|<2,�\��7X�~	4�����ͳ{�[:��Z���FjM���Xq�¯fE���=t����j��.t��)A H|�f�<��Gz.Ey;�����(�:Сq0"qj!8�ҿn1��˩��v��+UR��$\�H�: �܎D��RVn.��:�B�h�����:�=�!D_�;��m�iEGh%���.�8A@��1�P(��u��Y�X�lT!��7_/�vrZ�/�?j�aW��>q��\�x������U/6�/�-��W| ���x43X%���H�m N���?w~T $;��yF��o��&1,����KS�&�%dg_n�����z;%1a(�	f�O���u#���h�q=���4i��:���Յ�4DRZƛ�&&'Az�bA���)0����R�3\�ϜRL��p��@)�C<FU�����XH���[	x�X#�Z,�>z���-��y^���AY����������wh���j��+'N���"��i����8�RTD�f�-^��s�h	8/Mu@c�;�v����׿~�' ��}� �%J���i4ʴ������g֋� �IS��"̷H��H���O��?W��m}�4�&����;g]�kЏ�&���r�r�A2�FӨ:0 (��՝3�/�ǝ��Ԕ�m���xL�ɑ��(�:�s�ϝg�Zn'�锵9tQYN����kkߥ�թy�c@��p�?^�A��(+_r鏴�@�+R��h��e��. bZ|f�zqxrr2��I&��Yd(ɵԧ@Q���<�n�L$%<pzpf�����_5���"M�)؅�8�
?�k���Jf�	�;�6�����J��靿���1�ў|ù�ϝWB�{���)Ƭ�a�R{&A����W�����rH�����p�:wR,�̈́t1��=���5��3��hQ�H\n��TN��B#:�=�W/j�9��n�^{Q,30�����0!s]0��lҾ ��]�Q�U���O�Z �]����: �V&( Q��Ū���xX�en������y�0>2X
���v���	�*`t|w�[[[�i���TtP�n�@�&��@�CcJ����`������ �C����Ӎz˘kK�	�)�e�����j�u�`�`z'�L�|�u���"Y��f�P�4.$��%�C�3����z�� �/�:��7�L�v�|�Hga ��tĞ�Ƙ�+4��w\&v�g��uu �����:<�5�i�x��V7�J���#ߪ@VfzN��9l�b���w�/ģn��+�P���_�ŀjKk��C��`5������� )��Sk4�XQ�����ĝ�?�����KKK�B�'ˊ����^��ӓQ�\�����ҹrm6�;�E�T.��(�ѥF�
�%[�����Ɉc�?`c��>���0;��^Hd06�_�-c}�N�k4V�V�in.����T|syhvy(���+j{w��}�V�;�)�P&Q���J�k�;Jx(K�yxQ$E�Or����|��d�
��9	�N{��@2PJtf'���1���>���_G:���x�|�cs󠔴bQ��٪���ޅ�h �Y�������[Ȝ���K��5N�+��t�L���DW6������I�����>K��t�W�nT@)��f5�R��i�?�MXz�FFF�o)���;P<[����*m���z��o����p�X_���D�I.:��C�t�n��v�5w�G`�螜��h�y�]��{/ٛ���z���;��|!u-P ���KPS����
��k�RG�f��������b�?y֣Y��{��Y|~`׹�wA2�s��1�|��~4%%��ϟ׃���2���bR�R����m�Vq����+�.�ԳTVT0�ݗi�k��d�/uP����*��x8xL�[%hf>xe�Q��LO�%&�e����J�>n`����=%+��]�*����T"�������[`�cc��Aay�������5����j�Y��{,�Ył��n�́������>}�p����G�Z�
N&����^{�0�8��c,,�X�~H7׆����,�������*v��em˧"���ҲV�K�8S�Q������6��כ�8��ET%��(s��� ��Grjj��K~��${p�b����$L��������T�WB`_[۝���+-��$N�K�USUŹߥ a��}�}�?�n|�jd;Nm`��^�������X������kI�.�md��n���k�i��h��AUM��_��f�g�>�N�-J4lVa��<��[���<�@VAX�uD�ť��ŋ�K(��5oO��K6���67ݚ�	�Y�E			��+��`����>�}�25�GF,�,��]fE�N�YH8�d�A��¢(ȉ/����(|`֨�ob�RX�o�1���	a,JI�$�J��,�� ENz@�0 3p�z |22;7w2�A���mU��}����:�
��ZW\n)*
��"���EW�TN߫�ysqQq�-y��
�ձ�g�;��۷x�k|L�

��ׯ?�}t�,77��+e�/ .����]]� h(˗�!���/U�4���K߽s2�z��9�KK=VWW�߾5�5�`�-"����XL,,�e��Zce�C�"��}����&��� ���#������EEE�e��|ԦoRbc_�`͹��lQ"���ӮL��%B��#�h�o@g�`Q�D$]�ѝ:�Y����i!�ra.���/_~���9H�|O[c�g(ʰ���2�׿�k׮x#�5�D���bAk���x0����W��B޿��
��8'����o���8w�~��j/2�p��E��F����qt�;�������k�Ǣ����*ϥ�����&����˗oCZ��z؈kxGL.)��ջ������rx��h���8��=D��8I�xi��u�Ӥ��}w��b玢�6���[{��w/��w+��b�rͣ%�֭�?��<{�|dK������$��B���/K�_��2�jcն�.�*��D�-���.[�l�B����M^�������8BQ��f�f�E2&]�l��8�AE=$z��j-�x� �@J��x��M��R�� 82�����l��N�J�i�#��C� �|�Y�8�D�4m_�e������Ya������J+*�q&Z��]b޾=t�ȑ��X��< ��x�|	DW����-vzS�ؾ�DԵ[�;�d:Xa�=͓�,��(��VnR��2m~�K̘,*(К.�?��{�����j��܁�F$�f xY̠l��NT��`����y�F%Uy�]s{;�pw��W,ĭ��� �{SF\����J��:�c7��VBYJ�EY�w?0�������۹Y9MG�s"���z�
z,7�ikЏ�f���yV�0���=u%:Z$y�T��8ˉȦ�B��{�b�%������e�c=�w��.��,7��rH?�^����0���wF6t������G�c����#��@���Y}�W_R�Bu��\�k��!��M�]���_ ���2JCCCy�Ů�1/0�����n`"nZ���jo�_��\�d'���)��~2�0��ߨ����;���:�+��K1}��y��c_PM��v$����90��"��kI����|����F�bsU[;b�cV�i�$�L�&�mp�}ѝ̧����a̯��.O���.@3��=�Z�!�R]:t7�~���<B���|A���E�UUg%$zmh�s�c0|�@���ݐC����vPU��=4(�}�;�n���U6���=�>�C9��z�C~Um����,?�Ҿ�����%�^��:��Tz������0�ieټ��6RF�/���^�¬��D�5>�ٷq&�5k�� �M8f�L�f*Ԃ�r�;�l�6(�����Z�M���X�S������~FK^D	@�.�F3�G���h}
�Ȥ�`^]C�UUU�j�FP�{���΃�Ff���30�|��"k9��%��h�jtչ�~��������BB�r���Rl~���R^����'�2��R�c�<���J��������q�+�C�D%�!��%�>??�G}����O�Ja�!�o|}}!�1wON_D����
�sU����0���M��:l(�?��p@c�Fc�oV��Y�:t�8s��;���4јW �j`�su��\<N���^�.��
�j�G����x������U-u�	Jv��;L�1@���}���� ���'��?;zX9�?Yxfd̬f�Μ��j&�.d,4�Ρ/��4H����zT!\I%.&��������m�v����>�T���,��Z��.��.��"��ܐ����UR��܎��7�+�3Ȭ�W�G��_4������QNP<:�X�惿��Ȭ�{o��i6z�xq���{P�g���~�^��J��h��9>h|�~bb�O��r~�ޯ9��-d�+�(�F��I�q�+Z��)
��A!�m6L-Q�53�>W�%�����mE�%�����?WQY�����޶Z�;)�
Yw1	�Wtg)8�W���������h�w�3F��]�)�ޯ�!!����e5r��Zнo?x	*}Qr�@�J��� ���Ӗ�K�m�Z�O�Ϣ 	_�~�Fx�N�W=��	)!ܚ�Q72��<±��=�V��o���C��]d���;���6ONL�,�f���ŧ�?W&�=W��z��?�͒
ը��>��8Q=ܐ�D
;��DK�ٳg!*�Ԧ�d�l�(�ם��c,D!X
�a�a]3�Կ��MH��S_�c2�ĺˢ0#�"����߻�g��@�jkj��a<��8G�E5�+�A:e�C����q�w?��g�!|��-_�����)+*�իW�������
��	hb�q���<��m6�K-�t'�L���f�Ar4�p?�z�1�v��c,g�X��^!02�Z�C�PD��!0h;�~-+SB ��E�P$Q,Ƨ$>G.[J���={�Ov1y�|I��M�,��n��	�Io@��I�~5h���k+?3@@d�>{��>$��$��M����aw�S�\�C$���
j���B�����t}7x1΄���M%����M��'�\\^kl�'��fG7ۖ��>AP;�8��O�eG���y�����~���!~N��x�4z;@vZ���N����Wi�=M�J��@��eГ�/_�aa��_"��~7�&	T z8^��./�O6���$��'�簋-j��l���8��cu�*���U�����������ኂ���6]�G�P�A~Rq�Te=j&!?��"O�i")���'���޷]n�3�]Ů�L*�ȩ�+��ڙ3g`���?R�䮁�{;�K�7 �2���*f�}�r��~�d2��]���**��<&��0��m\Z3���Ǹl����t��PŤ5�va$���s�k�}~�o�c�k�<��z�W�z�Э�-�|���(�e�|���F���%�G��R�<.��3�3;ޠ
��%DF��ׯaJV�[�=r��"� ��W�@�A9%��wn�?崒ODo������PU�G�@@�(��hw]��X���iu �GQ�d�,,Zh��*聇P<�ƚt]f��>}:,p��ʪ ��**��<؊7�E�������S�/��~���1`�j�}1$��޽{:����w��N���?� ( ������"����.�CdX� k��MMM�Ӏ'#��qn?��!� >�?7?��Y٬$�;�&*���$��%����h_gG�s5P?��vphh��}S�|�G�}/�A )�������*~�����~�AJ��i++���sw���5ǣe#7�RV�Çǵ�V?�3���t/fs]P��0��?c>w��Z����+w�V�d�u��7p�ۆ��+��aa5�v�dP���1�KE��ߣ�=}l���&�!/S�I���%(K�)[���� -	H�nn�}!D�m����j��a&�L�YȨ�/�zs%zKS-^��u7�PH]\���υ�=�,�`��9ޭ�fK��72������q��7���dvT��'D�A��W�j�y�3Z�� �/ �0�f�}�ƌ�'ί�����*���h��QO�-*I x���k=�g99�l�P!�VF�P�������\��+��w^3C:Hr7΄�O� ��ׯ{��kGv:|��m����i���(&�����A��,y��uLZ����(.�E0 �.�>���f�'r�vCm��p��2�O!��� � �cQR�m��ݺu�"+���S���)ln��~*&�-An������ɽ�T��Vn`��~�osI�ܻ�q��gg �X�,�Kt
n�O�~@�.4�im\D�_��wk��Z	:"����h�{�؅��Lކ���qI��+���M+�Q��s��)�����M��G�n�Q��PA�4�j��$Go.$|�d�M���"z���P��	���������;a�?�����[	�ŧ�>޴v�膄���<vppXhw+�{vEA�$�ك�.��w�ܱ��Uٷu#�#�k�fı�W�_ � �9	����c�(ը�,��sFDDӻe�]�FA�ޯ8���&�$A^ꮺ���ZߖD;M)�
nQ�p��5�-%))������	�H.��v������'��^X\ZJ���puu=������	T��K�� �iiy�hD��/��y�*+*�99oXZZ��j׮=i�E�2�@��x�]WԵJ܊��^���FF�g5߁���ؗ�RƾT�g�`��B#͂�֒�jg�[|T[���g���F�����aM�T̬mL��)kh�������.����W�������/T�oul,�&ʽ]][�^=_!U}����� ���/_N�}�����Ec_Pna/wy�f=�}���x|Tr+�P7����jJ�J씇e�g)4�Etieuzk����Px�j��՞v���a�XD��%.-١_���T������}�dѣ�}En�c�ǋt��z044d`f�	��!t��P��N�X���Y�Ν��堭?���I))u6,�ԀJ�h�g<ƹq2���>�ڬ��e���N������S���hrj� ���v����+s#?�o�66�yy�߾}� �z�٨)��;"�5cF޽}��������6��`�lc�D��=���̳r(�ɑ�; +�ܡ�� �v^��}��1<���Ĵ��ZĦc���0�;9�#��������9>�3;''9%Encc���ӗ� �@)݁��RV����p�0-&w`~ea"%mbyv(>��3��ōiw�ݻw���#V_v��s�H�����s�Z&�J���_���[�%'de]jV��z_9�	��ɳ2�y�3�x���ϯ]$��?�bb2�nFt�����ďA{��Y0�5�Ӯ�Έ ���+�%h�m�Nc�sQ!���������~��K}�|��������׸���eӶ1 ������zz�---_@L$��1&[���i[��ޣ@�����yLh:����ȸ�樻�s�~��u#M�Vc�i�ZY��?��Z���zMH��I��{&�о߿~�	Ռ܇s�O����Ql�v��eko��j�������yyy�����2 �w�Rj�m�O/1'�͆�C@X�i�4`E����X������8��^?z^q�9�ʽ�����	b>s�l�oї��'s�k��?<�=~�H��>�E�������3� ��כ�:37w�}^�Ibu��_W��a���c����n��~.k3���h���5�Z�A�a���"j%�#�y��7�r�c�AV�B�ϐ�P���;�y��,U�5���ފ�UKP카[Ҵ�P��B��18�O{5�=��n+uz�߾��9�t��9h���W�������� X����>��]٦!K��}���h~B���[�)&�$�۟J��jk[[rN�t�qrrHd?]Y����o��뀡+�\|<Z)j3vpZ�Ou?����u�f���^��min�<�+(�W�(���L��@t�6���2��.uM���/����չ:^�ŉۋ��9�������I��
�3@���e��tu=��㔠��P��
�l~I�����5�Յf% ��
dp�͉��>�j ��/�Ek;R{�N�](�y�����)����Ц��Qhu��,P�Í�㵛U�K?Ky-���W��'��/=X�19&�y����9��7|e�lA@,�A���bJ� !���m~��A����h�
Z{z�Y�֟�pAQDDm9hjmXİp�s�����hQ��N��1PN|�t�xy��������$ �f� ��s#u���-��19��ͱ��gu�md�Su��y,ho,�(����[�Ν�71|���o��4v��|#u,� ��,����� 2=T���D���eV�	��?�W�o��6H��O���vs�q"��Tvt�����������c��t2���dC��D��+EUxX�F��������_[���^�s�B^gyx���+U`�.l���"b�3J?gk֓�f�s��c��9Աa�!�sܱ�;��%re����m=���U'�j������?Û`����Q*Ad� kX%�"�KD*��
dU 1�>�����������Fȭ,g�������u�� �c�~Ee��aH0b:-����Ύ6��X�k�ق�mNapq�`h��J�j�:.R���ɶo4�9��hsu��^{���oY���ľ�t�j�ާ'�� �9�;��I@b�-1�"i�)�	フ~���4�ƚ���,-�!�g�vt�JI��u%�Db�?L����u%�Tnm{m�4G�)C)S�M�̒Șʘ9dܝ�h�(S��9D�9*�g��Ӗ��?k�|���u��������~��Y�}wmm+��@ǔ� &�9{�]���˭̛�Mw��Z�W	�F/���<!X8֜�8�g�5���E-�r�;LO�� ���~�iB��M;�k1��G����i�l�}����KȖ�_W����=+-�=�{mN�$�m�YC\Y�F�B!?�u��NV�1p}K����qu���oVf�z��ʌC*�G�~0��1$�:A��{Rg@�$���8�zh��r�&<���ep0D�����Ȼ�n��)0ȵ�W��<v��[jֈ$zӶ0=tkn\�{�M�����&a9Xj*͂|����b��a��ЀEC�����J_�C?\�����+@U�]G�pI���h�y���Mq�}����*������Y�utq}H�z��j�)Q��5�&�	$i���,���MT���.8Vׇ�ʴ�=u)�~4��m�FB���N��3���9V��f���uuOG��c���	�U{�����c\�� vv�������bh(��.���Oo�߷/ğ=�
 �i�����_|�?�+(������?�P����iC����)^g!Qv��&�~:'�8ȶ	�Q	�50��|�8t���<m��6Z���ю���.���䱗SnyFk��Rr���pOj��p�%"""��'�s����>kkh|4tF
`ܑ�tӤ��g=�\��r�#5!b��tR1˃(�{����1f���F �o�F�<~��"8X����3,��e����ח��y��	�2���7���7o��_�~ӁW�@�� f[��i'X�\d�2(t�8�y�ʕpЇ���ݪ�n��e�$�͛]��H {��B�I
�o��W�\-��B��A�DY*��z#>� mxZ9�����[@<�`���#��v��4��np��AͫWߌ\F��2�/č��壱����D�ق�|�
���5a�.@b����m�_{�t�>�>γ6�ֱf@B\ɏ?>:ڜlii��y_!��7�7*z+GHkC^�f�	�vJ#pe�$�b �,
"&"'��x�r�wO��=k���$~�nfyR�{�r�!�6K0�('�gdl�)u��9)&�4�1ccZ@_�h6��x�J|�r=�t����C�sP �޽�����ٳ��1��H����C��b8Q�y�B%%�L��q"I%o��a]����ִ��0�([arm�K�W�+KMU�����iC;�"w�hJΏ#��˹Js!�p�0�����W�c/j�8"D%%�6F�����:C�{���\ݿ��t���9����1�������>6_��G � ���3�f-�0c�G@P�<�&f��k�t��\��ֶ���@R��_�}	r�ʕm�Nt/Xe��
��>�r~X;��Yb���5�?�#dt%�y��۷O`�^��V����h����2.�D����jrsR��s
ؐ[�}���I��!3�Pi/�b{���^�z�p�G`=�A���8���Y ���mD�T�v`�K4d��@��Z�_�^�::c���<�]h��.���OD�]Td@�L�\����z�
��`� ��9��!�E���Jg�/�C�sE��T;v��.�-�� ��qs������cX���m��5����['���VjδhT��r���B�� :�??�������J�󄦥e�d��!cN|�C�[�n�y
�QE����ד�^ \�N:m�k\��E/�x��.��2;�:;$���!�imD��j3ʲ�sΤ/ݷ'�UMM�uqvL��mGH��������^��l׻��g�_Q���؋�P��ҷ1؝�R���<�<b���I��ZZ�z ���o��E.��_�&g\W�6�3���o���٨�D�dNLIQ�-^�O'������� !د���5�ٰ�.���H���^(ZH�	��i���]`˾/~y�q��������Q��[N9d�h������_��������k�e�*
�z��E3>VB��Kz��*� ���,_TUU)+�os��&��غ.���1��(���ݻ��}�F�1����#���k[�q�����`��x����0�ql�+O��ǧ����_���Ɗm�S Q��{�Z��i�	�s�ؖo�G���8���X�p]�#x�Leƻ�� ?�=���SnEF�@O�y��͛7��_Y��]<UQYA��Ն����A,���M?��˝�}��"���9��Φ::��1O�>@k'
j�{ho�v]L8 �OD�_�		I��R�oݰ����M]M- *eSOO�Zl�0�k9�����d��؉��Ւ���"kih<Ղ$�i���-n��Yf�ܴnֿ?��]���s1!`縠� 儅�n˺X��)�nr���/
�/�:Y99�PU��Y��� |wV����0��t����Jjj8��1X�a��'':sԆj���N���Ȑ������c ffBG�Nsl��=X]n���ޟ�%�����O��9;��m}��SƢ	P�`���\\\�n�IP�*X�sO~�p����
*�Pѿ��>"?_�sq$�]r��(b���pS+���Ħ�W��1duWMu�_��Y,��b�#]���Z�ϊC<����-�����
�=N%���ІM����Mk��'�t7c��{�������zp�JG������3�q��mt*��� �@�?_��������yk���c��bR�� �KO�Yt�>
.mc1;�Z�_Iڟ������*�������݀�h��ċ�z�X�.���}k��aB1<cd�%S�a��w߂E�:��y��qϤgiP"L޻C+�����JI��p�8RQ������:3�Xr<�Fwwl�ݮT_��7�]��.?Y�g��ri�h||,��C�`n߾���$����˖'h���+�5����; @�<�J���66SKٲn�jOf�����wR����B1_�i�o��<2c�w��:���?�U�	H#��%-�yǁ���n�0����ǽ�8��8��8��=2q�z^l�I�Ӟ={@cs�96:
2.¨E�$p��o��I��' �u¶��#x��+ⷮv��8o�rb�((�acC6OT�蟞;5����u�*�Hbq�!��a�ΫܟA;O�HIԊ�W��`_��2�Y�xj�h_�<&[#��`��'�;yx���7��{m�F��������|L���2wƨ*�4����0Y�l ��ޮ��`�	ӱ���-����4x.:��A�gJ~6B���(�?�e����Ѡ:i'/�NQ�ql`����ܻ�#�w��#�{�[) ]s�="%=���e�ǎi� � *��+3c�,��h��!����)!//t�{�:(�:F�ڸ��G7�{���;���������43�.h'Р1y�CAOs���C�e,��t����оu+7� n.՞� �r�UG����&:Dڠ�c����g�e�Y���ǭk"e�`!ٔ����������׾nf��G�}����jͤ��O::~����8(,�I(��ک��)����`"}e�t�� eNA��"�߅�����Hn^G��S2�k���\�����lp��Y�C�8Q&�|�c(�?##������; ߁����Z5(W�gyyKh{T�j��i���,�W�{8�
'�G��`ƪ �׺�=6�d2�L�)���M������bWCͅR�h�T`ш��g� `���WE��<��l���g!�A�#��	Y�!�Z����ޑ#���={���Q$�8W�K < ��DE���!@����*���z.�w��d�q���|�䔫����.�x\[Ay��=��F�[9��Cb�yp1�hM���\E�4���i�w&>/ X�U�h���ʂ��2�ol�q�q[QVV6.�'7����B}0g+p�7��A�B]N5*I��x��%���j峈�Lv0��ɴ*�|�7&P_c�/U�J�LW֪.Qo�b�L2�"1/O�GK[�E�A�in�&��?��m���@�y�)ۅ�=#��)6}�`|
�a��wיִ���۸�:�7P[[����/�r��ߍ3U��ǲ�Çioa�b^^C
���QQ���um���v��)�?511�+<333<�j�
|7U��r��J�)��k��,���N;��eEE��}�;,�[�|*�WV�0���A
z�j�f�	L� �,��ٖ/++�:88��<(!�*&��bZG��9EOOO�����S��}{&��v?I�VVY7;�4�D翘�����J���i�;J�ϟ,�^��M�}|{~��1,�a��Of�������mڲ%�%O�����g�ZU���F����@�o��{����_)����}B��Y�ش$�Wm�����o����\Y�v��j�r�HM1@n��3�o�q�a�g��������&M����5�\;�S������FFF��6z���_��9��>b>�b$Q������eJ�?�qk����@"@��f��j���8{��������l���Q>|�H�'�����_z	U������իz:��������5��kjoO��qI��jv:�uT"h�溺h.�ʾ)�^J%�W�ԋ� 6��Q��022߹���h��HH�8�
Xx���<u٫���1�9T����}*<%��k*U�>dd�����,���#�1�ߏ����c��M`�p	+��a��uBh��xp�>F�y������s���Kq�fq�0��#����> Z:���O�[�l=��w����W����ٷ	�I1���v�~��}��ߏƗ��߿f�:�����|)�rԶ	&��ir�dƩ/_}{v�~=���+q@{��X]�,�^n{-.�1;�=��b$EQ~�!˂���z��ffj�6��2�5~�"�`���ݓ�������p9n�q�+)���֭kz�&�{�I��E��v���ߜ}�i^���nvv|	n�]�#�K�_�.�\l�.�/%%3f���&��d���/�^�▓��}|yP���%�
��M :�htџG>5F1@s���M�#x�����q�;��45�}�*�_nI��u�ӟ�|�ӧˇ+�f�ѣ���]o�II���V�	��T�g��\���L���yܐ�b>�{��s�g`��l�o�ј}�L����;�|~��8�	( $�IOOO�_�$cH**Z�p?~	�O�7:|x�#��g�/q4����LY���ggg�!;�.fkv�L���vv����<N����.|���C�o�@	����i�ϩ�Y����/�
�?�b�Ok�fY�T��;59�Յ�!E�AT�%���9�_�(��Ŗ�b��0�cμN�I]���-C~��(nPľ�{�� �qw8����ѳұ�Q ���+`������Z�麼rXM�jv���M3�^���7��#��9WX�H� Թ��>�xO{���2?�j����Q�� 
�XC��tz�>�0 �J�W6���&��,�0�.��hu��۷/�,�Y���/�Q;&��	U�K����WMM���%%&�/LA�çm���R���@Z��Z|��|;�U� ۦ��g| ��w����4⨁W��{�.�M��2(?m������,_'�䦻�O?~|4�d9%���y|&��qoȋF��A�r�p!߾��4������Tm]]ݶx�"�������w���}���Xk�XV�a��D��p+�ؐ34����h��@��i�ן@5�wg1�PQ���J*�B����s�	�!�0<�<f�	j���g�Z
��T�xk�ML8c���Ђ���3ާ�[����)��������?��S�����c�~�HmN֡�~Z�o���0�dgP��B:�#�&{� ���`.P��C}rȻ����뭟�� �q��������bn�A��k��i�2���!˪UY��A���Ԕ^ƵG��/���1�ƛ1�S��ȏ� ��c�����◬��=Zjro񃱠�������q��%%ͥ���;�����f-A��,����Գy�<��TP��P�M;2%����4)�h.���"�f@�YGC��J{�JJY!���o {چ�r�F";�G�|6B�	�y)o[o�p�elHHH���%�w��u�����:���DyO�[�r�;�?���CB�t_�?L��+����HV�W�����X�֓�'q<��y��n��Gp0��M�$�ۂ�o��de6(
�h��!��ٴ��U������<( c��g�,Mӗ^�!s:k�(�����ìv����i�W;hm��נ�ҀS��o���μx���0@������I)�"o]���*=��s	��q�6c����KM�����`�p���6]�^B;�us3�����U�[�(�}���-�`�<�8�͞��"�tHt�	�5�� �����8�5��5�(-MMџ��\Ǫ��������9|RZ `�n+��2�@�j��FZ�{��j��Y�P�� y�o�(z4N:v40-&�4-$<�ti�ٱ��]�n�ڳj��H̙��z<�16�dr��?����<ڀ�?��~mf�j�m�&�����s��L��h5��?#	~�R�?��\��\!����9ִ��ӣ������O&>��e�K��?\O�,hhlT��!"6���щ�����6�wc�6�#sss� ���"��t���Wǎ�����q{/�ӶF`��I�z��؂6�,d��f���'�v�Ǽ�YR��?o�'�C����a�MwD-ql���s�1#��D��ܦ?�0[�!��$Ѐ#���b�X��D#yǡ�L��.=̓5�����8~�H��FJ�����W!ľ<�щ.��"�N�^�[Yl-���u�IhG����n��'�f��Z?2����g�,5����F���tL:'y~J�������zs�K�#�b��t�B�W]�m�;�j���+�����ԟٯ�D}DO�_�[�5N�!Ҷb�=� ��k�8Л���c����uL>���� i����n���Y�C҅�J�:~T�!eѸ�jҳ�9u��7�\\(�<l�CP���
����wj�DO��r��C������$�x���;�����?��υ���xl�b�7�ϣ�F�h��),��j�����6���ұ`�P�m���<�X[�Û|����i�܆�h����o��'�c�!mV_�Փ�����s��_�a~٫�1�;�a{h(m�H��<���9��V�
�v���-T�T�<S��M͹�_�6�g�����+��yw�����?�xD5ƻ�����d�ȩ���W���]�_R�z��}6��'97<:B��aLɛ���kZ(�5�UV�I���E�V-M�L�r��&8Εmy��D��)�I[v�ͳ/��o�@�Q>�.��@W͝��Ȧ��G�o[�b?�ܒ�@4��R �����@❋{g��U�f�����mݽ{��,��O��^���|��i�ks�XP�Y��Jn/�̢���H�$0��j�ɾ &���=�!ݏ�u������T*�g�P��WK3#�k[��-���
Km�]\��6;'������9���G�������@�V����E�XO\�B,�Dnc���^�,��Lذ��#%��}��9�c�W�'i?��8VB�_��Ϥ$%���$�M��qǺ����S��>�u��Ґd+i�n��2�~wiJj��"�4�VOG��_n���ܚYT����|��N��Pd�z�ڧ��#F��F�--��v"��e��!n-���5 �;���o���:R��M+7mm��,Np+*�	��K|H�nRRC�rgI,�a���I�>���������i���X����	5��}��ښj�Ŀ^Pi
���IuY^���]�E���Е�5rw��C��=߭t���v�O� �=�/�fCM���7� �{Z�@�*�7�(2G�p�W�H�,�@(���8� ��"�W��"�c�I��\j^)�]�qdf��^%�� �����R�u���[J��t.�4u��g�x��`8\(����.n����0=���g_O����K�\��/x�.C0�I9���[888�3a���z��'Pf�_@bF��/��-,�������������������d��^X�2jg!
a�%Ȳ�)�`3� `FN�gs��+�mm`17����+���&�P~�=Z܌���yw�-e�m���07��.��� ��F��y�1�q,���+fvq�8��P'�3�/Z..Oz�p�#��$:dӻ�0=��S���rt/1X��2�n���ϟP�j`r��d.��B�t�eڃ��T�fF���03��m�&䬊�B���׶s�6��{�*�z�7���_���������^��/l��pp�^ض����%'+�~{ D����<������i���ylV9���l 9';#�9���&��<����:F�Ǥ��]����Y��m�_l\�$�XU�&�:bQH�5X�C�a�_3��Jb��Ґ<� !������2hmm��^%iv(�r��䤃��K��~
���v�Š(>�\����r������&$�m{]�=��	5�U`����,���8�-�!��s��G"�P/�j�Du�Q����P<�<��
�(�-ǘ��%ʹ0?�w`���H���
B��c3%J�2� U�T�Gp#|�Ĥ��J���s�*p��%<\5��2:lB��?�C�+fzFF��ҴxE�o�J����p�(T �ȵ+�4\�D�3��ӀМ�����i� 8�gF�qg�r+�D���J��N`�Y�*:$�Ub۰��ťK�ޘ�R�v]zu_H(�
�y����K�ԑ�K �؞=N;I��SqeP��^�x�]�r&q�:����a'����
�}��b�.�� 8��ƿ�RD%��-�H��5`A�x�<�ev�y��c��.�lz�c9j��gY� �a��z���}�z^+��7ӒJ+%��r �o�� ��y�c{P�V.��,PVqYYY�ૣ,(̥o�xm����g���0��B���1]3���L��fo"�sa!�0�l�a�m;i�u�B�3�@�k]_��Z~t~���'�����mP�_�1�^�o{��i��"j�������MI� ��~*KoN����?����yP����^��~�9��8qb�PY5�-��1ͼ���:������@��������
�) _eU���P*��`9�d�j�Z�]. ����.��&Y�_f��y�0D���;�bI�N�j���F5�{�e�O}0茨y/j�=E��D�Ӫ<���EC�M�q�����p�lʓG�֗��v۷����cy<�ꏠk@ȈC��	Gǣ�
�0�S@��i����t�il������۸bv�dAݎ}[�(A���N+K8P�������z�㣨���J��� y��{�M@�#�mPIN�
�!m'4,�#�Z77�}�I�4r�T�(�.\��u��N��9ƃ52>�9���"ُ�Ta,��k�m��q���p+���
������uR�h�c���DZ����:�߲�O�����s}L_'�������l�Ph4|^&��-�"�|�Z~7�S^V��N��Q��%`��L�"̪��=���-n��ʧ#Jy�폅hwmJEh-F�͈�BN_FG-�{rcL�e��'��7uW��jeex(}���"���:�P�m�����*B��X��p�߸!���z���Թ�՛�ք�jW2����#��z� _`	ByҞ�#��_/�G⵴��`ﹿʈjA�?�Q��990){dw��G��@��-��r��"|�Y���&�D3*��2�i�V�r�2#�E�S(��f���޼�Qn��ZǨ�r����O��v�c��Ǐ��)V0�A6��9?AP�R&">� e�f���O�0i-&�B�d%#��.GL�*���d{����;�N<à�+��6�@*Z���z�}�|0}IWW��B��e�Y`�ͥ����{H�Ay��c����~�u����̈S9�U(�&��Y�%6y��hk��c��'�a@��wk��T[�s_��8���ہ�M̶�.j����<�f Ujr�С3�L�MZj�II�d���((���W��| �p�=�w���4�l��t�v����[̤��Ny�"��筻��
��P��Ʉ�x�j�i���y�fd��h�j�_����-�������ӛ�xrӱ/8��r@]��k�����!�%"��[�a���}��mH��'O�+A��G��!L��j�����Xnq���P�Q���r#����ՠXvq�=��v�Mk[��`�SDLf�n૭8������_�A�"E�i�e� �����S�]}m���.�����_���֣����(wr�M��Z��.,�,���V��(~Eh����չ9g�[�0E�ZA�&�&�� ����\�q�*%ڶ/;S�:���|������B:B�"$Y�V�u�|����hK��#��@�J�6=(�Y��)�~�
���U�tX�����2&�$�W�w�m�z ��O{�j M\�U�qD� �7������ad�UG��XT�Q���V�/�najʇ�%0y~#��ʟ೪9�(Sł�ʰ,��o�O�=wN��� a�,�Vu�����"�NQҏ%�-��U
��qǇ%��n���풐Z��.X����qT�����]F��B�I	�JR�#1��R�	C�a;,M����3�/c�`ҧ!T���U�p�N��������F&T���<C.�C
a�hvD�BF��AR�;T��&��t�8s3��3�(��Sv ���'>wƽ�?���?��=1���pc�T��
����
�]Kz������P� a2��\�E�Lܠ���"�vް�2ȵ�+�E���G1�+�I�M���j	���ԁi��h�H\'��$>`�\c�&$��+�� r�di\s�
$�%�&T�c1�8�=��|'\���"	��r��h�[�g���B��d���� ������5��B��(��Nd�>޳�P*WUJM�S���8z�"$���D�RZ$�^;rwP�d$_sf�Pz��_����+�h@�����`���H]`����tu	��n����9���X�z����^Q@o���Bk��5OSN&6Ja�t�J�!�"�j�} �Iy�xШ�+dnB�������ѕ+X����9`8�����t�0�#. J�C.%T�u����$}��En��-3nEW�
�<h��2�jKqN#��N ^5���IÆ{��ts�;7>���o��5ۘ#�aH��з9=^2p� ����T��������oin!��=�@��ς���;]A���J���$�zN�@��#��?H�e"�Y���J3">x1��.�ٶpJ���A��N�PB9�U����~0�S	��Ǳ'�Ob$�X@���vd,��?K��Kj`�$��QV��^�۬%���u��=k�&>�"���Y��r+��A�m�~����s5��>�.vOz��eU�
n � ��^�u�5?�%	R Kd����~��C)��+9Oi��a6?��|0���aV��ߟ`ǻ�s��e�L@Η��F@�A-9�5��ұ�g�� lӺ��v�.�5�H�#��\d�R�?j����ߚ��X���i	Z�Q�/��H�AQ���}��%�P��{Y�P�<N����}�N��P���
M��ޢ*���l���
����P�CD%]��w����;g�J���c*�zO��^*c]��ó����1�'��R�����fԔt�����j}i��~�V�h��v
�,�.L���P��mɠVC��~}`��Y����]�+���� ���ٌ��>���<���0��]ӵ�<\��FQ�>��<h�ف�q�y�d��l1�|}m�\��)��o/,TB��_4�����ן@|2��o�Ou��U�L~�<������w)�E��L����5���v:;��T�������P�W^ZZ�QI���a��ԗ��?Q��]�l�nTZ8P�%����w/�!�Q�"�6�!ī�d��eS|J����=���Fb3��vq�h�^G@o�����B�dݩ����S�$�ʿ�j���z���w�h�Tls4�v
�$%�W-3)DwBigAո[I��)B�t�ҳ��"击�Á��-$�o�͗y.0����-���FvZk�i>����ҧb���	(�,Y���q���[���j�g�d�j5�8�uE����A���_'P5�ڈ<���Z���]%��Q��\�5��.�d��.=��t�� �)Z[H��˔F������S�K�����O0���6H��l}��� ���Ṇ"g�<��_��f�"�0����u��u?к���W�4���͛7�V���ҡO�n�f�/�J:i�:w�(9.�L/��I�U�1��m��,$Y�N�N�0 �Lq�zc[��Og[�9Ze��ۅ�:���Zo ���idrz�3En�5�~m��x7�.V���@���~�}>2�^��������a
U7��{�,d�1��_к�����AN�ʃOJ�z�t��f'�fgrW�;�uRQۘ��5���Y��O�颍1�w���2B���6ep/V�����`F<ҿ��Yb$Pw��#�:6+���;i��G�THi�ݻw��C��]������{@E���b�onQPD(Z]џ�<����W�D�]�d;����}�ΰ���yQ2.��t�$�Ā�I.񒅑=$)[�m�|�O�Ъ5�Ό)�]4��J�T"4���A����:c'���^����|g�.X~n�5���^�����!
�mH�����d�����.��n�)))ץ�N�q��pz���eQu�����T'>8$"�=��`�7���s��@urZ�e�D��p꼙���@�Z�g�)3|��e�S_8�I��$伉�� 5��J���q�bB�@5#����?����ŀ� ͗܃�s�;Th�\�i�]�@���{R�(�jaa!���\9��/�?h2�cS�^�m��,��w�|�VA��\z�n��g�hޡڨ �.�(�K,�A�P��[����"<��r4/~�п�a�й=��rEOOi�ƍ��c����%��e��8��޴�Q�0��M}����-�xmpp����H���8&9�M�@d��^��~�ʕ��x+��;��|Ua%��E0Z�Xo��������Ӻh���_����X�3l���Sz01�Xq�FsqfՋQ��T��T&@�Cfum����z|��(''=�X�����E�F$�L��~��Sjg��td���Ś'��=�dZ�lh������0��G�}�.�#x��+�IEE�3i�G�m��Q�����.��A.=���J��Z!O��%Q�BGC� $�����;��|�4obbo8���1���d����EE��	�CVv����s �wI��ʊ�B��Mv�E�����Ԗ���ш�)�W=p�x��>���(Z���r�j�V�lz�?V����ړ������$X|�ZU9x����6c�8)S��>/����O�Y�Hvv���_�o����Õ&7�������� ���p�1��4�Z/<y�j��U�֋��~Z>y]_2��X�dr�=-�9�\Nz�bt���$`E�I��$ߔw��q���L6��\d�;�9�Zge���>Ph�>�yB	MJ�kh��
r[��X�,Op�c�������H�mj(++�_Y��'�O
U�`���j}ocUzf�L�wˬ�u ���SW�6�:�~��.3y@�t:�=�HL� �Q��l�%���2.^�`#�:&\Q��n� �Z�z!X�s�uv��)_L3 ���*es���|x� j��H^%Q��~������Ր�[�x��⬲���e$P���/������q� ��݈��h���;K_����$H#�tO�9�·�{����-�7t�##�^u��id���e�����u%|VU�z�4!Hy�3ql����D{��??�"c�8���+S�e�|-�6ݺݗ��#1�9�!J��`���ڒ{4�����e'foǈZU�r㛺M�^kh'Rײ���`���o�:��SA���"T����(&���6�0C�v��^6*�4�A�8;
!��+�Ȃ��EE���fi=�u��Ց8�_;�>;�� ���I�wO󖧩))82o����q$tt[Vy��6�j!����C6���_��H	�aDƀ���5�y,�7�9������ �p�	gwր���k(� C�Ҫ:�	>�����w�g� ����C�?�c��>#�v��S:"n��D����[����i(к����� M%���,��.G�r����~�Ct����{�s�}b��{i��� 9�����=@G�qgL%���8[��Z��Ov��t�߀H���kE��Y>:j��S���5��2oWn�LI��&��KP� �	��@B^!��L�l,Y%W-���(Tl.}QĶV��^�	By�I���l-.y��TI��TlpA�����m�ޭY���?h?��k�:���Yƃ��V�#R	�B�ﺓ�7�>a2�c�e��bD���!��w-�v`F����T���=,�!:Y,F��f��_��?6���,,�]U���6�W}�f�8/��f�d���;����#\��"|��g�64�a�e뤻2��w���ĉ��s�����tD4TY��-�� Tz`"�N-Q�����7�\�zwp[/�M��Gl�޻��s��'ӆi�\ 7/Gf��8'ڕ���o6���g�/����E��=ۈ)�:dI�����	���U�^w�o����S���{,���+ʺøזJ�����#���x*6�'��I��#�f��UM,�tO�{D��,�n�_6��J���B}ĩ�8�fI[	��9|$kԎ���n��&�������d��".{���BfS��澘D������A��L�d�$�B����D��������{��Z����v��QmX%���0:I����`Yuk��Zg��}�)RD�"+�D����+�X�ù��w�	���N]4S �l�kssK�g�,%V TTL���P���J�r��[XեR'J�Ò�U?2�+w�Ȩg��3ãh᥿�[��}���N2�`}�0�F���j��Ω��,o�#��yiU�r�#�Wv��r�.��V�2��E37�sb�ܞh���NMJfʒ������9�g�Nu��[�!����yĒ�b3D��mP�^iኳy���	�[��}��[�-�IO �(ߦ��E�x���%�o�8;$Gl����m��x2mh�	8��5e*�d��O���j@?KQ�u��+w,���D����ؒ��3l�0w��͘�#�v�A��lռ+��NQ�4P��х�BC��\L�n��<�X�h�-�B�2�ə�iK�&�̡n���zԤ ��qUF@�cGze�Y��\��Q�P0gt�É��k[`��o7�~ߔ�YO�,���֡�8���)�ԝ4ˤ��"d,���h�}�,��h���\��OA��:�]k�5�=x�<�m���2�jk����-��� mco/&}jbi?7"u�����)�c�y�$`=�Kۆ�˝��4hE�I�k�������E�u�)��QL�(�D��s@��Wcȏ�}�yGiW��^���K+	e��X?|�J	T���M�^xj���Y �}A)[@���Z����܈n���c�&��>�e���Ə84�[h��+i�8ȈHΉVT��{��o��\*D{�6���W֟x�w�
c���+�#	���:� A	x�AoS����?���ֶǢq���cˈ�޷[����*[���(\���~��D�rX2]3��j�_�����@΀ ���ݰ�\x6˸���&.�Iy�.�s������pǛ��B~����Յ���V�t� �3�]�\��c�5z�n"x���i�q=9�	���Ä�W�4BB��ʍ�R�WƖ�ҩ���&���P=�f'�������}�6�u"�uJy��_ �F&M�Tf�$�tÇ �}3()g��3��ɡ�@/S�`�B���r=3���������0C�����	����e���`�������Ç�*&��]G���ׯ��.��	�Q��nƌ��t-�D�X�3>�7�m�z_qu�t�1w���u���(�4�gh?<:�|��Ln')�8�$_q�>t�W\�).p�k&�f����4�p��SMlP�_����II�8x�x��D;k��9�!
���'9闸��t�ҁyx8�Wa�`�q�뎴��A�槚�fߘ6����E���<I4L�zJ|5ܓՀ/���4�(��`�y�A��e�ݦ�d3���
,��@p_3"��j373s'f-(�1��r�	�O���;t]$ ;Q)n	WZ�A����Z3�@n"�i����
K�DN��7�bYyN����p��t���	�paĉ�+��b+fjsu��Q�O6�å.�Z3�9 R�V�2��5.O�1�c��"�OMn�?P!���3J��r�M*v��R�܋��R0c��d�m�d�G�\}ur�w9%t �j�����FY�l�DT]J��v��B�'���?mEw<���@L�3=�A�g˫*l���,V.H*��P�
�����j6IIJ�#����<Ϸ#������T^��� �n�>Spp����@M�������q?����k)�.��p�$�:*��<������~�&݇V�ř��!"G��\
�a�1��&td�(ۙ
ɝ x���D3���������Jx��8����ώ�(m��n�r��{k�8ѽ]�6������m,78��%���	����g횿!�D�vQT��0L��
���������Nȕ���'Q~�8��P�5-�7�ݾ��L��q����;A忖o��`|;��X�]�d1������Cڡ�;d��YLE�ns~���=M��_{�f�8���9��C�����+A,kks^N�@�Q���*p�L��VE O�����M/�<���$�q�儲��2s���J&i��9s��ǏH�����ަ���%OD}�_K/�b-a��Uw�Vk��|w�C��双<��ek��}�(B���(DKP�����H7$S�#�QԮ�ɍA�R�\�ِsVa!'Wo)M=ך}�Kgmk+a�~v'�ή��KZ��"\%�_�����=-�{pȭ��\��E^��'s�ւv3\��W���'	}�`e�S*�(�\�w)=x�:��&F~��7R�����*�5Ù-�b��U֞7�����*�@��/q�-��fW�F�*=�8�y8;3��}K�u��Jziةx0��ɢ�hՓ�'�/i��2 �F;I�%n��!T�;B�R�b��b��[k�c="���%����C�|�hQ��}AsS=MNֈAN�F�6���Y���C.Y�v	X�K5~�bo�#��4l�j+?��M�e��9��ӽ���7!� ���S· �'�/��ڭ0m����eQ'�dd���go��{�v���?l����j�Xģ.�6��3b�8+m|��� N� 5;
��]�|��0m���D����n��1 �&��`s�f��xYiY݅��cp���)몮���*��.�?�bs7E8�a��Z�f%�_G�e�!c�w�r���a&j�ج��-ZW��JR�����k�Z���w[���&%:������X�䣭��y�9���~����xT���N-��=�Wq�8|�8=���� ~4u0/.|(�U��m�'�ѱ����9e�I���͉Fh8 *;'gȹ ���1ɺ�s4s�Q~����w?����׃G�U���nEy]B�d�Hw���'f���[F�ٵv��M���q~��cK���,��#�֫���{o�9��(O@��a��\F[SZH�hG��L���ۺ������7��A�O!F<B�5����ͅ���K#OR��Ԧ�E6�1�8���M�f9�N+;��,^r��yE_���K��H�Kd��F��G�ck�ff��ʺkeW՛L&�M��9��|]:������)>�wO�c�;��H�;��Ql.R͍_� ���U|��f�0jy�lȁ��j��������Z�p��B�)���l�����n^`��/O� m6L�j��Ǝ��J߱(~��`qI�q�����?]Ľ����Q54L����S3�nU�y������0�{�Z�������7����	(�e�"�^���O�'Ri[Vk�W<n��y��䤃������P[����X+�;G��Gg� C��w��_�yNJJJ멻���z@��̦Ix�"�P��y�"s+��K�ܶ4��۬�bcc���M{trPP�m�����جՍ����[����|8�hl��F��;�q����'�@\�m����ӻ2a��.L!DG���uWA'_��I~SӘ��pߨ��&�h�4\�G!���k���|h��8_�[G�@�����������������pU���dev��=�g���1*t8#=�٬��+�u��f�io��es���G���Gz�.v}�P�No�m��DΦk d��%���M\�x"��H�x$G{@��8�O�;�2�/E�?��}b:gD�h}3?������%�Tn��/*%q*M�J!"�T�y���yf��%9%�3��d��IȰ��,�!�2������ߵ��:�\��]���׻���G�X|�w�5�)'QW��f���E�H$ҁ3��%Q�+���i�H��U�aξ�>�t�Gi]ў#��q��Z,�A���׶�!Y��wa�N�nN�$7�
���� ��@��|.�p/;�WL�,�ʳ��[\kֺ�"��U;y"�x.s�w\r=�9��
al�
���f::7_v���:ж'Qoz����E������ߢ���L��c���7	1��[��Hƀ~f�����1��b&�5�F�b��[���ԫ[��~�MfN�k�z���r���~<b����>znڞ<�a�wޟUnK�G��z��NHcG���>����ZY�$D׋]������"`0�g��Q�1���?q5ky5���pBZ��m;��������`6=߾�mqi1Em��L�g�	��H��n�,
Tm�7Vˌ6���~�h�ػ�K$e֬W��O�aԖ�y �#LMU���	/��#�v1�}�Dc�R�K�R���`����u�o(5^n��70@�y�&;+����;o��&�l�;�H-��`X��9���_����!��f�2ҳ{�얃r@���K�p�05q�Ƶi�KL,z!�ff��Z�I=�� (e�)�
�g���*�G�"����?]YVvg���w+$(�yÖjQ��s���ϯ��� o��P�	�$��+x�d������མlX�`g���ȯ͖�"5�O��i��������X�.
�+w���$������Tx�3K��~+��k~4m�{�nݕ��d�V$�o��T�Mj��� _��-r@'���Nwd�!�g�+ x���t�tu�WWZ��n�mq����^��O���0su�T����9�rS/d3C���-�]�}.�|��(���c`�Жe�l������ҵ�&H8��j�I��whh≈݄�l���Z����	}a�N�mp�|�?�j��[�6�k���;�����Aa$�q������-s=�_6��Ol���־����։�&3,^>O���d�#��Ȇ�f-y�x�:����Iu� ��vm�;7�[B^1��cHO�a�L�NoWJS��B sّ��o�ţ:6X`A\��Ξ|@H�=A�ى�����XSU����Qk��
ePw2���e������œ#*��#9�X��ݣ� 3�>M���$"��t�J��C�\�uVC��\D��N=zc�}��x�����T��R��B�� � �a,�����t�Zk���\��H�%Re:�F���T���C��P�#_no�����F�C��)eI<���P��%>��m��F��� ���t/v}D~��'4+<�,@ �g�<&�@�������L�8�Tz�ǐ@��R�����eqX������9æV5S�kW��}boO�#�[�@����t���)��B&}��r���y���P��|f�@#k��+�
����|��A�9`���A�dꅛ3a�(&[T�R��ټ:���I�3��q�b�L
��t��▦�z
vcm��2V�����ׇ��E�L�� ������ �pOA ;>}����ܝ� ��@�>�z�Y�=�<LW{1杚�yA���F����u9I�/�4�=(��w�K�Ķq�;��y[T\�ӻ9i�}�8��U}�e�.L1v�\�j�mv�m�k]�x�C�4�zK������e��ɔb�c���&(�Ş�� ���9�X��)��X��c�G�sЬ����f����Ŕ-Pw�O*,��E�$�q�KS������eD+&&��,�yRlz��}?{4�A(�H�MEU"Ǒ���ϯ��D�����Vm��|4���ki��F��+��zl�j,y��O�_���0���\]��l��Ѐ�6	���U��_#�2�̔&��lo�#uV�$�J<G�a��]]]�U>r��Q`��=	I�_J�4vV�:lo�l��[�z�����!�����^6�(z�$1w����m��ꟹ_#.�k�1�Kg�ԕ�H۵w�c.J�]ϸ�oEqP�ᓶ+}溫�����O
gϩ����;�=�[�����a���VC��yvs+g��sV����V$*8�T���y��)sD+s�ĺ��z�I�����('�@p�~�� fÿ&þda\�⹱ٯ����^酟<Tpb~)-V:���&�1,���Y�wK��9�s���v���Zl(�ȩ�ڳ���N�u�W庑���櫂a!+;[%��D5"�|:�7Þ2�W�xm�s�,0�T�uQQ|qC�6_���	\��V��&���`A�	�J�9O�4fC�k֊<�b�n�u�䇹��Q7�j'��u��5if�UU��pU�'S[E%�*�.��3�����;�𭸕�V��S�ɏi�[����9/R����\E�*K����Z�fw���v���0�9��v�y��T���;5t/����8&Z@���¬l{���Z��{�7o�'���`X S|r�)�z6'����q��-�gu�.��%\�_��DZJ��n�r�*��S{�jE�1�|�z��T��TȼI;��Z�>���M�ye���=I,��Coww�L#Z�d[�S��-���P������υ<ݽ%�L�3X`�0f� ��L�����Y�h�D��>�am��޽�V�j�#����m�{S�l���W�����Yo��JL>�|v!t�fj�]T��`��f��s��EP���_=��j��Z�^�c/�u�xr^��K�\⸭/�Y{����RX�?2oӚ,�O��<��z��SŲ�ĩrFb��1����4���P���FlϹ�V�;�4���R��)K��ރ��@�x$�k�[]zh��I/���x9'�]H&�4���׻�Ч@�%9�V@�S�n*L�5��~���X"���I��n�$X�=�J����%�|y!������x�ח��D�im�Y[+�,v'+
Lv�+�)!>,u`�WY����f�[�v{
̅Y3�{�O)$ߐ[9��]	%�U���NmB75��R=�3~��$����j�+O�1c�M����A�m�|+ri���Ni�1���W�<M_8<޻�E(<M6���(��6M����?��+�2@�jD+f��)F�t��f�<�� h:D�(Q���[oUN��U�	巄��'���OЅ���
ݔ��0���(2G���+��EIQn\�5��� $)�Kc�Y�:W���\�S��nzf���X��޾�������b{2�	4����������A�>�+��涬xr�}�����@]���g���q��	���4�W�K�v�*��"�p1>���|݋&�����,V�F���%y����=���jj��ǆ�`�(_��H�����߫�'�x=+��%����C�ُ&v�k�L�9�}�X_�_VV�v��a�1�(�.��:����UJ�p{�o���_,߀��d���\[�j��<�PM�#�.,"«��Dc�첑sU�Y�LV2����x�5=+�A7������ ���c�wc�wSs����0ޖO���,~����1��N�Ƀ� y�]�5�W�LiY1S@���~[|�I6�n����Ǯ�0d���
RA���Y���H�\;�����o�Jϐ1*3�S�_�;53P��M]���HeBh��5n�x .����}��/�$�5s.Iի��>�c�{7)��^B�II����z���Mʱ�:&�����嚖����í!P��Q���O����:�M�[vl�"�bK2��^7�Drpp@8�@`M���F��ŕ���+��i��BT+Yq��ׅ1�)C�<�ݫe��e�O�a�ϟ�w�k��V8R]V�h4�r����M�,�A�b�"2��h[��{V���5��)H��Mp�xb|��L��ɧ������wpC��4��|r!�d�-��[2[�����3*jj^}7����J����.W������ac� ��ձ�?뎔S��9�F66�|]��� ����_���Y#PA���xD|�$�l���b�;,N˰����pW�4��u<�N����@�b�Y$�ԯam~����{�(�J��NDB����/d�o��^ ����-v��%�>�X�ק����X�ľ�Rŕ��jL����t�\�tD�\��\g�e��̉�K��=��ZMN�,y�1��б��:�M����F%���9a��/�+��L��V�ݡ���Ce�g��χ�<��sde��L/�7'=���I֨��V�WJ�!�)�.�x��[���q'B B��}��Ñ�K%Px�U7o����y��a�۽c�2)���M4���I���ӭ_�&|_�j�/��x9��T����J}m�)fuL���|FO�e����I�����|GC��`�������3����ن9���Xgރ�ʡ�J|�[�ϖ=i^A{��tus+f�7n| '�X��͝71�T��g􃹺�ʬ�+Fl�?ɷeb
�p��p�D�XE_^���sx��,&:u +%�1�i}�'�va�2e�(0�OmmO���Ğ�hx��!�X�6���[���W1''�G�طg���K�� NYr�`�T*�d'��E�f�5���7�x��$vT=�Sٿ$ؒ'ύ���w����y T$�b�{�"K�v�N:������ijfa2�b���Ҭ���g��PY�Kz|�l��O��ѣK.f:��'z���n߿mA>�:��a_��[e��6 |��!�	K&?}�i,o��nή8�SC�N^ד.@�Zy]蔑���� ���h�1��%��#Fڷ6�Ub��/pE4X8l���1q���*��,���ǖ���o��G3+6��ǖ�b{B�Iԩ���ʱi�<V�m@���s�M���2u��/�|�@�K�VP��HO�mT� ��d_/�fe����FA�=��ݠ���x>��|'�?�d>Z۠;}�4g��
��1L�Ub'�qBpm]}"���XU�X�/C@A�8�5T+hP�ͭk5� {�Z'(0�����+<��2���b?�ig<c��k��و;�a�Py�/�o�����>Xc�ŝoV3�ꆗG�Gf�a�� z����ܜWO��fw�<L�} MmP�D�#����r�\��O�^� Ps/�0�ws��F�(@q�,~�:�� ��Ӳ�+ݼ
��Bp�&���PAW�]�\�g�5�y�"X-��b��(�*>���	II9=k�'�F~u#J��a��9P���b>��q�i����*����2z!2�	g��5�`S��SLV'�&�2M�� (��>�N�ϯ��nM��a@jB kQї�eĩ��cb����%�b�&d��<���r.�)��NrLc��:Ӿ��k˷�=τ��^뿕����`xE�9�Y��E�
�SކI�Q&3N?�W��5}��oݓ׬�o�ʡ{��d����{y�G\-���1�h�j�^��YM.ϛF/�lnn��ҬC�Ȋ���ԙ�%_��'�By/��f�����w�n��@o,��X#���K{�A����3��[m�p���"F�#5 ��i� (�u\%����@��b��0��*�� !��3��B�kK�b�F�u��6Bv��������L��y���&�J�b�'�4�x3�&1ȋ!R�L��<��?�#�9;}Aa:+b�2A� �h�=��d���V~t����+�Bi��Z���Rv9��{�q���"���.Tl����6��ᢁ��}+ ���)�u|�7�чG�_u���@�v��ľ�ۚ��3Kjzgt�(�.���	{��1_"�n�z�v��C)���_����d���,{1�ut�Di�g�n������3��/k<*WPao���T�'�e�Ko��r��q��
��-�Bz�5���HI@eX̳jڽ���������b�������yݣN 6:��6�#i��O����f�Pa���\b=����[y\/��,��6�C� ���x��$�x�,,gqԘyrnW���B���љC�\��+yx<�<��0m�bx���o7{]��\���j}�X������� �LE���a���;�[�U��f��J�U�(<����
/�@ M��������4�]���lK���߀}��=B��U�ˤ]����dڏ=,~��b���*�owx���>��z�A�f~�^���n-�����O�*��/a�e_RM�g�.�YW��	������'I���7BН����=�o;�]�rܞ[��6� �1���k
�I������Qy���� |Y9[�$�L,�U~99�W{;�Er`�_������:1d�#Vm����#��~���� <H)l����.�><���?��m'���*�c��PF&&-��	��.寮��
��dZ��&�,�z��5�Z&̈����OW�Lu�bX�tJ+9�c>�/H.��AD�����{z*l�"���<����G�f�f��a>�(?r ��t����s���Q??��t_#X�����0����;�H)}x��������(,.���aQ��a	��m@�X\���+SW�{�����Tr��Un�vz��u�+} OJ}͚
;�D�u����*@0>W�F���1Y���.	���9�wVB^Rb.,�44Fqv���~���֯"3���oP��RG���U|�l��_�:����G@�](W��4̅���֨�9�Ձ4���dSG��>MO;�����p)�G=z��s���ئw� ��-��M��Wg��z70��^�8��]����jd���1��V{er�bq=_�0��4�ۡ	
��n�X%t��3�]&��W��H̎�T+y��T2V�稰�H�b�-dݱL��۷���x�wt��H������>�ȡ�s�a�Y*�@�Tb���a5�ad2��l�6_���D�f�mt�j���m��xǿ8WA��7x��H�AAC\6��+���4�Ӗ������� �u��Mni�oU�<�h�oy�DD-QT^�ņ��&s
t<���E��w��"�����Q�@�lB�6D��eM�.��?�C��wAI�׏ `Ҏ�]g t�FG_ʌ��OxJvv#���mr��ᄄA��w�e !��1ߐ�D��etr/�=Y���~�3�x�	�޽{����P&���EN�s�-	|��9|uu�ݚ��t|���y�n�u���������I/�¡���B�*�?�O���5���Q_cgg���RH���[�Ę���o�L��v�c��p�i���o��=l���̧�ڍ)ˤ�Sj�L���%�ޒ%`�ܬ��ܘ�����)��]ucw{9����}N^J+8��]��2`��Jل�cxO�����	Z�η4@\A�$�R��ճ揺�+�+3}zJ�o~wy%�$,"b���	�a���nD�7c�����>���o�!�;��T�|�kR�[����+�Ln�/>}�D^|��&�����6����y'BWA�o�Ǽ���`!���z�M&ߓ�}v�e���9[�1r6`�t����=f?c2o��]�u�{巾,&¼��}��b����v���|]H�-*�h��e@�������b{":�^HA����A��1lb�D��\"�3Z5.�ק��J�%����5�HMy�n�'h!���oGk��nG�K@�v���6-�K�̺��X_d�ٍ��N1hŠ� "s���G�
�x��5t�TQ��m� � �����uO�~Y�����(�`��R�6GT���+��Ǔ�=������S�6�j�K��߃��p���䰚T�:Wg��4k�{�^�*S=������n�a�-B����~������&s�fn���ؒ�9�(;�����K�=�h�b����!��E�a��ĉ"��&��6O�'���ݵة��8�P�*����������������V�]�Zo|�A���¦M��T�]�W�@G#P^�������ӨG�(d�ʺQ��Ea��'PaQ���N���Y=hn^��[�^��V���EA�΃OC@6�;0��]���&�>:��W��OԼ��Zz��������s��{� �&�ر��������z�\F���w��؄`����T�%M�Ɣ�;�]��W
��m����o��g��$�u8��H�QuI4�$����F
P��f�[�H���ӓb�&�9���?zb`Db�(���f�@!�˴�ó2Z���@Wi�h`/'2ڔ������GC;I��HM�H��$`塀d��\�WD4:��ff)訲���y徭
�9!3i�b͜8��Y :��.w�&ɥ�jn�f��8H����7%�E��l�<�եX�'����^=�	T�EG�ғS�Ƒ�����M�,�����b
h��T�--bǏ>���nl�[)�]c~A��O�ȣ�i���f�J.��q�~T�%]����MKax��S,������=�b����Y��cTh�Šy�m�)$#�0��A��O����i���/Z���މ���f�@��,�hs������24��c�-�,J�'&��g��=��&�.��s��_F�}GH��P��y���\�e��^��6�a�7��qV�[47�R�c�Ձd]������#����WO��-�����,�f)�Y���Ն������c�N�XC�&\.-������V�w-.
�n/<�~�a��ya����5DOҿ(�D~.y���hi����D�xXt&S�@6T[M�W�0\>>|�G���ІQ�߯�Z��HQ`U����j���$ꞽ�˛I�%�	�͙�jc>kȫ	�rc��!;�?����.R�@�6��GSc�lD�we�0�O;�!}xx8k�ko�O�E�a�Pؑ��\�nhe�G���Lg�\�����^�Kw�
lC=J�Z�#,9��W(������鿀R���=���g��dG:��|
c���9
�q�G�CE@6D���l��E?o�3s�7D���]d�P܌ t�c�A!�~�Y�zl���n�\D��t��j�߽�C�b&2:}jRVU]���7�.זb�m09�e�_C\SX?�ǅt���l��L��>l�_g�ȉ����-=yo}i=�#a������&z��VߡGf�+��\J�y�0`$��<���F������a�γߠ"�O-b^�_ԣ�%ڦ��&2"���D<RL��	mq7|a�h�r��w�c���}���i{�L��T ��t�02F�yTD''�S`^S2am�s+�)�:9�Bi(�!���M�a��v�#r�t��ߑ�
�~���N����J4�9c.�P=g�A��:E�?[�X��	 ��[Z���V���T��22����L�ݴ��ʥ�OT���/�8���8�2;F΢a)���%---k���V�1_�R,����a�aN*��s������g��ŝ���N��56����vC��he��|ʚ%�'L�����?�\1s� .�l��v�M/ّ�)�
'��2��8��^w���uS����z��ncn.�_��u���}�U���L�>�����ק��Q��$hr�G�)�[Ǥ��\FPoSh�"{b�Q�=�Fȴ��ߺ'�
s�r@���8rs�2ay�������|MHݮ9LB�/V�;Z-�)�u��ۿ+�o�ņ�Hfk*)�dK3����������Ŋ֭Ɏk���t,RI���l��|�-·65_�k�q66N�8�^T6����K�~���Nh:�ʬ�^[[K�P�>�,5c����B����b�p���e��~��ǟ6���r��֧�!�_@���^IJ���;�@�,�,F�=�%&������p� ��O��+�J�;�/��])V���3��?�A�� ����!U��뤬���P?}�,��O�-[-`1���0��������;R�� �}�)R�ל�Z��g���]�5�m��o	��'J��%��k��͓j=EC��%;�����\mn��Q�S�{W�+�(��z�C��?�)>R�,���Q�4�X�1P	��ÉSp/	�����6�e�f��U���9�am���G��� jZ�oo��If:��(�������bAv� P&��'CBKB��=��ڟj�����D�i�C�t�������c=а�o���~����)ڐ�У�2P3x:�_`�A��s�3?I�?���sD��g:��������;�h��������8������uy��)r��jᏆ�g��Kkd����R!"��m����9Ip�Q�L�ى����O�>�������i�˱���
��������'�(���_�w*EM;���1�����y���������X�B�����ńԂ�.�(~�%�J��.����[om*^$�y��1�V^�V	���槝���~���ј@�#.f:�NO��A�hս{���)���y�@����$.A|N6¶ٺ�e�>�̾��vQ���G��d������om�ru֖���͉#�t�R�0�$���y�1YD����!�&P�l���ˍ�U��>��W�(7F�ND{n�� +k=@�����\n��G�&l==��L�bQ� K�����C��mj��lKn�H] Y9n)x�D]�j*d�h�ߍ�5�
4�Vt����D��+8&����fZ�@�&V]mi W��i�b� q��v��J�r�n�{�[�x��i��F�r�ɘ�Wrk�������z���cX#�=eY���m�Em�L�䛯�>������'^�G)d�~�&s�%N�lK��:� M�B��M�拸W�i��g+�d�+����}��L�c�y�����I��V��wfΒ (Q���g�*�})Y1�����௉���W��_@_���4��«;R�]s͐�!���ow�g�j���@��#�c�֋��[��)^Rg�*�K�Ѯ.f��X(��+7��t�}���u�hu���{��+�����\ȓoR���b� �;������M!�?QKI�>fz�����d*l������Ǥ�P�#J�#�Y�. ���Oڶ����W����c��ff�:��w�X��7YYE����Wrb�2��\�-0�A[����P������=�#A��I�F4d�s��ޫ�TX�4Dk���"I�{�'��%�ݟW7��DS`���I@4�/��m`�QF�L}f��\k/��zX�+1ۘ���ge՗&X�Ao�V��=��&���c�F1�,���>�,/����@@��R�c�v��,ߴ���j���+�^�����/&$%y��A"������)Z|0��kH���U�S>!�<J@i��=N	���>���w�gbO�e���Ǐ�yU/$e1��3��G3����W�;�%𐱏+;od+�j��ʥ��_�D��F�_��s���CBBď�ڎ�Y�ډ���v9W�^�~�{�}I�� ���[��9�R�{�� �ѸheKs�$(�Iӣn�q7��w��~� �0����K�9D�XHm�BΡ8ħ|ד��RP�(�ź䆑�B˦�Ꙛ;Qci@�������w�A:?'�����9�66��e���x�a&���c�@rž�8&��ʡ�V��f��y$J<-�C�j���6��6�U��0����E4���$%�L����ˤXk+�@v��`�5Bae0�
�]`XGV�<��ӝ��,�_#����X��y�*�l7�/���W*[����(D$X�&�����}�FT5����AE/Uπ�[3-�:,K��@��R��������{f��]��0�������T.{1Z��d�|�+�U��A1����i���S�J�~i�������� I���6�}������ͬfO�^��	�ɺņ&b��$c�nta�n7��r�
f�Ԍ�O�?]s�������ge?����J��ɿeG��G16͞5w�ӑ�[��V}A�� ��W�P�o��g�ֿwst�@�p�6�,poV.@E�@�?�wn{s�J؞��A�ᓄ�h�D4j֫&��B��-���H�R�H6�Q��t�di���ּsŐ��;=�W����ўZ"�|1j8��֢�`G��M��[�#i�CP������B�j��E��n���9!X�8�x۱̸��WU��9�rZ�GV9]v�&���*�^r�#סG�k�;u�.�����q��0�ZZ��v�ا>�Ok+�٨���$w��B�GzٜM�>�e����WG�)_v���� �qŞ��gA�;�JT�s�`D�ϩ�4�3~��C%�N�{ �X�����
L*�,�����+�9X�ʝ���ydZC���W�y��/�m�A���a=[3��h�a~�fNs�TX��}A�{������4�� �Sչn�gad�q WFM��dV��W�I�1G�[_���{&dF���)�w&y�P���Nc��k�cK��0i�v�6��6]�/ �#0��j�>�[�=on��a������������?�&�6�]��e�=6;��8�8�3�j�=gʤ����u���)`k-��e��`&�Ҷ��	�?.��۠�.���	���ג(J��]����b���w�]�/Z��fiP�������[�W���[�c<,��wU��C����)y]SG.ᵹ�6^l�Ԟ��u���h�ȩ�B�����3�Z�v(U	j;�V_���m�l�'�4��	�����d4��'�vv�O|b�K$���X2��&z�e|a#�����˿m
�������qy*�"�|�!�Pk�h惾����j6�<�G�O9��h35��'�$D�r�e��W&�HW6*�+s־h��^T�Rم>5OT��W�S$;��W֋�`�|�*�~3��/Ĩ��y&_��\C[ʺ3��_�'�xp�D/�
:�����I,r4z����\�@  @�i�`qx�8�<�%Gh�qm�@�~� $B�|�������w� �q�}��R?ݪ�R�ٳ[�2����P|È�Ѩ�q���rz�k��}p<�7��Y�⸾<�6M���uo|���z	HTKs3Wl���9,�C!u���"*l�J�0ox�h�<ݾ<Ӌε���g�Z���ӈ��$Z�N`.�-|�4�v��䡽1��%���(�q�VU`Y5�-θ��g��dR� ��v�����E)�<���Ap����7+x�t��]	,8&�1�IV(;;&#��@yvQ�<������:�\0{=[7���$0�$���=�^�߷~��L�F��M�0Q`.�~&q�����)R��c2չ^^?����J5Rw�E��p�0���!":��7͇b.�����td��)P�P�oWKb�APix�j�9Ԏ�; �g)���{�⨴�ȧ0L�c���J��o��c�T���M�����_yNK3�����J^��m�^d��%�(�\�:�P'4Vi-x �B[d.�ͷ���ޝ���g)Qb�����ȉ3a��=��X��TD��H�}/���z�Z���	����t���8V,|���-�,�}r�<�Ǚ�b%��g�
5�q��iTS�UO���
L,���G	�JEE����\.��ef��L2�Ķ��� �	�������kx��E��\�E�z�W��ZF]�&�Ug|�r)��azz:�����@�~'<V132(�R������T��w��h'م�H�%R�y�5�2�z- �XU�Rmm �tu���y�H�ݦfu,�c�o��)��ؓ�.�ƪ����j�=��W��i)��&e�E��~������q-��ȅ�T�k&������V=��2�g���h�ʣ�E��!h���.X�����t�n@��_��C�z���`�Z�]a�"�c�/�˔�0��\ڐK1������ �zjj �0	�e�i���),53��p逷R��];j?��0Kܘ3���1�_������+brFA�C��g9��}�������\4��y�/��8�����9�r�BG#H�a�;��a��d%!� �%��B����0�
�dG�� �g���F���;�D���=���0 �q��g��9���xX�a�Wi^}�X�XСgo��*���[o�x��jP��� jV�2%���R^^��66�PQU��	�qtށ��-��Q��N���-R�iS�_뿽��u��}|ۘ���9���3n�ag0�`( kK$�B\0��M^�o���[���Ȁ���w���rim:+I���80����3	�]�F��eDq���؏Z��7�+3̷�uK����z�I��0Ķ��`a1�W���\Ϯŀmq0�L"�F��˟o�K�1��]J������L��ш��$/;�'O�(�D�����[�������Kx�B��q�w *~[�����������1FBBB�%���+>����`����ɑ�Kݨ�oĥ�2��/���]�""H��/���%@�(r�8@Oo�4������ޞj�����j}2h�>��\�������J���Mڢ!��Νo	��������>��� ߖ�\O(ԋ��)Qj2���P�v�J�S��������XϽ����=�9Z�8�l�25��N���z�/.�:����� ����"�y���33�F�o�K~^���O�n���g�������?mh����7}�Hg��ɾX�v��@M�{��n ɞ�ϻ�UrnbnkvN9�������{�	�b�P���uGt%ڷ�$h�F�J2�)���9�I۹�i"��	��U%�I� �i��{�]�}��x�:�3�e`a�"ؓWD�����E���r}�1����0�,�DtP�-w�2ʖ��k�0�v	�DG]"Ia�m���X~�*![X$=m�&���c{�,6TA�Ѱ����)�'�t,�-��$}k�D ���: N����� �n=����u1��b�=�Z܍	M�]zkkn{ wB:�����2��l���M��ܾ��^�Ԙy�{�.������`Ƥs��Q���_u�X����J��3�8�ó��V=W���?ژ�����h�Y7d���QI`��3 t�|���>��䨠��E��4a�k���Z�Pi�|�񯓙�����'�$�-* �P�@_�Zϲb���Hx��Ԯ��޾��K�%J���Yebo��^���P��.=��D�����e����"�V֙�R���ͬ���N�7dSTO-U�M�G'���H8�6��3��!��HD�J,y3�ߟ�d+��ߖ:y]�򟵎G7�jsG'���8�3�IԮ5Y�����"Ʈ���!qpʓڈ��Wȣ�(�ؑv%�ȃ��?h�N
��y6���^���9KD3bk���I�'.]7ꆢJ�{�p&G��s���LLF�^�ƺ|�Z|��l�c,�l!��ƞb��%o��ݩ
d�W�i귤Cg�f�3Y{�
5��<��v�\#���-K;3�Հ�?d�{��fIOe��	] �JW�.'��#ɱ��忒�3����bx�Ȥ	d��CP��꾦\£��u�c;@���R��鹏�&�Q��@��5����:Bz\�n�=y)V�����k�J]�Ko���t	�X ����q��v���C�?�x��Q�I�
]Q 0G��N��7����� �j�l�׊���@���A�Ϧ?�z��N���wu5%X.
Q��\
G��X���/������J~����1�<���j��b�G&H��f���[T<���&#��]u���>��Mf{ϖ�O�8�C%��g�|Ʈ �N%6H����B��e�j��%p�'�;�_�"d)Q�D���~4�b�{g�}��V�z���I_���ݔ�F%�萪 ��<!�"P^Aa)�m������I�7P}z�ŧ�U+��e_ض�(l6�l�N
z3��2�8W�]���ڷ��N����S�A]N�aC�����ۛ+K��̸�y�d�̅�����8J�b�QE0��Y���c�m�8�p!��?��7+@�
@$d)]f:���\�j��'����BI��#�n���-�@�c��٪�����!����Y�*�k�㨌�9�� e!��� ��$D��HW�Gh��/j�ĖSM��`;���uR�m����������o^0|��(�R�{k�A[�ÇQ�E;���/LkMf[�+�f	II&m>M����4��7tcI�F湎�r�( ������[ڗ��u�B+���o"��F����;!3u�1_�lͶ��h0�wFĄ��{s����f�?����b�6L�
��\���|*j���-�gg�ws���	jK@�mq8���s��y�Is�~
����;1�4�F�����1ߘ��܄Z��fK�zX�u���}�k��s�W�f�˔���k���#+�YPJ��D�Ψ���̑%X-�fee�7�����s�(��]҈�""u(P���b#d֮4n��}+ f	�Z��2 V����:��z�v��w�S�j��bۆl,��������8" ��BE��]��6��2���d�[��!��l��������jW�\Ac�}�����[�	�Q7�K[�K�f���}�]Vj����%�������oQ_�`�i�z�k]�빍횯���U)��<t���oi�鯸��jD���,���^hpފ#I&��st�u3%t�s���>����<ٽ���'�9���z�ǡ��"_�������Y;p��8W6%���2��]�U�\� Es7�>��ƆoK�Ei��pJ�%=-�2(Nͻw�&����������:�^�n��t0*22���ѱ1nNN��/����/<�be'�������7Yv���{LiQ���K7��v��[�'D�E����ͫ�F��Թ4�2d�.ʊ�{��h=Aq�Zw�nnnT�utus+*UTTƗ��H�Q�)��I���\Q������P�ȴ�������!�gׯ������]Lk�����,;XZ[)\��p)U��e�(��1D=�4�\	�`�֖vE��,'��E�*Z���+ׂ�J�r�md��uA���а�۷WccV���o��y|��?{�4 �mmm�|��ne�U��]tRR~�I��k��ZN~>�ǘ�P�^<�.9�~��#\���6�����\I�Q�st>	_S@4Hʑz�oIUC����4t��2?���֞�5\���#>~���>*��_---�WY�TUR�|�hΉ��8qLW7FPP�a������H��}g(Ac\;�0��<�Ӄh��k�zm�)�c�=��~|I�. �Xv����e�~��|�V�����[_N�fbbj5�--)��̼#Q���u\B������%>�
.^^����l�/�[+c�����8���b�
�4��r�.o��h��5Dά�=��9Ӗ�Kf:::�Crp{��NGC#����
8~��C�HAU�{���}i�T�����WTHq�񩺺�*^�.�4GR�������b�+��m�ӧ�/_����W3��������sH��&��{8���Ϝ��=%�Y�o�Gض���߄��Ƿ���Z_�^�f1M�4*��hynwa윀@�&&S�����76s��*,ԄyI���RO[O/��'��M������� �n�[?�X5%������}���UM%7ec�L)�o��8nx��bH*?�N��Uf�;A�mf@M���+	���'X��2�c�S�4[(�;˦��c�5��K��EI�9w���`�v�=�2��G�x:kI�r��f���t��^�����m1����U\z�����2�E,�xㆸNAvVV�Z�E�Ԕ����u�Ý�c�)x&��Q*�`�ڪ\�Y�{����F{��`mj�Б�=Z�W^��M�]���C�uVz�]dUd����� �0��b�SDxii	,)Q|l��Vuq�S���_�[S��5۝�
��'�Q?���H����қ�"8�ȝ���Ra����ۛs��$�_q.b�Ǔ}Tњ�Ѿ�)��,�\�i�RY����?P��f	�� Z5�3�h�/\�c.�` ����_����r��<������������-*`�烍FA�C����R��D\=m�JhG�Gm�ҺM�y�.+�ϟ;g98���W;?�LS��9��`�ѻ;�]+�'��Ҷ1�����Z��W��H�D��N|�TJ�xQB>L�7�A	�g��>�=�>P�S��8]X(�>��~���th^��s2��-j얮�f$��yJJ��K�� ���:E"�����K�~�w􍵨�l��ͨk�7��۷/�����-7�V}e`�Z�-��{B�J¥���DS( ޴J[[{1lPe|�����発I�՟����lf��}sf5fQ��o��|	2�~a��[�O�|�f���Pa������To�Hs��������=�u�Cz6'��˽�R�����a�N�T��ض��
�%%��<��pu}��g��qyd)�6���DZ\�u��	�!	�YY&ٴ0����z���ޝo��a���{�x*��\)J��HR�#�(�NHV%;�̤̌�(�쑑Y�QB٣�}p22��뺏w��_��~��<����}���z���u���~�܏U�
<�~���bw}+�WI���K�����k�&�J]���a*��J�Lo�ں������uhhH���]~�7�錿�~�0�~��*��tq�L�,��sp�Nh�3�;Ժ�I�o���Xo?������i�d9��w�O�w��C]���I��r:5����Jɵu�Y���G�^LHH`�p�AE�X)q�Lw��"}75�����<���oki���xЦaT�Hj��6k�x�؅�4����l��Ǐͪ���?���N2h����������5�𣁘�N��n���[Q�0�R�D���vG��
'SK�vC�D��rb��G�@����e���L,��j��]B�>@��詨��-�g]t�3̡���L��ϑ	��a<���F��R��m�ߊ�S��B{fZ�T����k46G��"B���42�|MW7���X"�_W�"�7�屏kK���V)L%x:L��=-�h��uNT�e#�Y]X�MU�x�q�kUZ���B�XCd��A�U;�U�R����5�IQ.�~|�5�V�0Q_eq3	������x���ե���uP�rb��ղznˣ�0^�Sn�ףһ��-���GP����@�04���ђ��n�q�ңD��q��i^]VPP ���tuц�Xi�tK�D�kh�-x3�dd4��@H�c�
��*xmbIɹ����eVf��CC���{�t��Mf'��'��W�ퟟ�\�U�!m�k�ɍ���7��(����"v�&l4���Ag�~m��=���,���V>}ןQ�O��AQ�|^�N������L �&SR�88�qr{D$��
]�$j��a�b�)ʷ�N�eML���ж=^��,p���e�8��� �u�͞��2��ܬ��N���E���)-��� M��-ҮY��r�@+VD7qj*tdTg�_rgf>�g��oA�t��P��9)Ci���g����$�ۀi�0'3����$&~�׉�122k�[ip,ۻ�m�@K���G+�Z:5HD�'5�o$8�?��������y�a�����z1�Ps�ɓ';���=Sj�INӅ$�e|�Z�]��#��T?H����6c'̴��ph.f����$�!XvXBBϱ�)������R�;Χ8� E-F��j�3�u���pb�>���ø!�Yk"���ԂQ��k*� j
���;;��0��BIa2++kZ��ǋ�zo
mI)&�QjO>�:I��F%��YGł�x����@��S〞�������� �ݟ��r��#� �����nz�}ظQ��Ƥ�{��W��� ��G0G�GN��Z!l�P������:!!U �ڡ��w�D[��<���B��"Z���p3�X��Uv!@���� ��v����9){}��^I�><MY"شʹ�����W��CJ��	Kk��]�M�ɹ&���Q��Ϡl������#��G������a@h��jp�B�/���/��s���k�-6������D��'��-���i���t���������
�e��?c�r��&��D���g�7P~�%����q��ZK�su�#p��p��$���#,�5��.����TG�,&�E��� �*���#�&� +�	��O���}yQ��;uapZr>��s@O�pG��bIO�+����;և<����� ������z)��x;Zi���,��r ����c^&:m93jzb��y�uC�)iZ�D.���'����$������u��aT�i�� ��_�3�ۿr,�Z�K�對��n�>��o�nys:�^�&����� D���	Yz�[*v;~|�W�5�N�M���]52J��GoL��S��/O���'''��������?��� �vU;EL*<���>����h!�oE ����9�����Uj���QW�f��n�W(k&�ʲ�>����8�0�*�Z+[�Q����h|�(��}���8¤(�+���bE�3�{JWə�}��C0D"x��qP��3�+�X5�u<��(B���Ղ�*"N�8]�p�2F��m�T���j���k��Avp�	���p�*)�0ࡦ���g�sH��/78*�����~O��� 啱o�����2{��v�ס��`����i5m�@�v��މ1��ɩ����a��ɗC�
��~�� D����A��W�~T������߉�y99B���{�|����q�$��q��2ݞ��1��^T�B��]C��W�2�э'd��'</.Y�՝���EDn��`��t�LX������篜���K�[X,~:h��sn�$ܹ����	�Hd��Q�
���n#��a��;�.���<�a����p�����d��c(*��2���0t=���%���6��Zh.�W��'.ލ��ٞ������B.�X0Fy��7$����ZP�`a���Lf�NZ�����I������_:����e��rE�p�B���WJ�c##�`���>l�����]�<�E�Y����2�L-r[��?1up|�#]�ɩ��� ������p۶, ZI�;%��fhx8�0f��SU���[�w���8L��=s��Ѓ���H/y�'���-v�S77W/��@����R �U���M�	M�R�`R�2���qb>�D{��/�!�jF��Y�dD'��i�����QԴR�u��Eֳw_�v)�7-�W���C/���9�
m�����ݨ��QD�[plPH�1��y ���D�y����R��`�<�u� 7�����S,k&���~"�.�G>=������goaa�#���w'��z�;�><i!���	0�����,Q�Xy_Y3C������=�\;C��?)]��cc��8�!�h��)���� ��m�_Y������%BQIU9B��z��z�����z�g�\E;�:k_	2����uP�u����F�]�ίuu-F�z��'X菝9ӊ��VW�s_ �VQ(�9V����󞗞�솛�zKJ�"�6f�lf߳��8P章�#�ʛ�:�$z-&Z�����(���ՊN�/2>�������r\Q��7		|||�0~-�k��9�����ǵv��_r�g�4&g�i�������g��]%��)�p���^nEUMMͶN�V�=�X�TDQ^5��%J�H|��]��ٞ	+�߱�[Tn�v�Vu�[\넬�����qE����z~����?gT���.�#J�ײ>�$�1oOS�ZPu`��E럐C%J��.��-"҉��5ت"5�vMdM.���mU�Ȑ.�+�o��pEI)����p������p������yyy%gL\Rd-�I����k��&pIj:�3K�Ԍ�]�V����!�����b��s�;O	�� �vpiD�1$2����"�+_��'N9�5ee�k�v��S32���3\@EM\�;�a�"?�#�>{����gO�S��W�M��"8�Y���֡����F>0./�[����=5��
������_����R�do|^30�-�m��$��0a�8��s��P^111sr!�g	���tEڛ�9�Z�R޾}�����۷�:�7v+7-��5�$�d�<$��餭`
O�������Yv�y,�Z�sj	I�򕳔ȼ�R��j�޴��H�Ȇ�������X���h��ƚw��i�v��Ɋi�����	s�D��]HӖ]%�,�I��a=���o߾����կ����⡃���h�{A�toq|^���q�#kpn	������Y�`��A��M�z<V:��Xyt��JJJ���7ᩣ��}�Q�^�G9|�YCM,�>]��rTW1�!�ԴSu�XE	7�u��/������v갮ek���vi�m\�_��:g�j}��Ζ���"�'�j(((\�x*{�+�L8Ӣ=w膞��ZA���T��������gir�i��GKa�##��Q%���i݊~�O������sx�O������P��"�M�׮^���b���DG�]��˝��S]	]]7���A#,@#�|����ӣ��\�����R`0jZ��S�1��G_�Et0Q���@�zvW����	qqG�CBl�v8}�	��Ѵt�|TE�P�}�KB�Tw~x���:o�OXXU����>���0�����&�y<��d^��$0��֌�i	
��kK�Z�e4`j�޴�Y���lR6R{$mq�1_��\xbE;�5�nֿ�[���c"QMԗy�Q�/���]��L�w<i��qXԚВK:K	�Ǒ��\��i�8�S,���{o�;���o8���[��s�NCqO��W M�^��ߪ��ne�a�Ŏ*I�����s��ؼF���o߂��'z9l�D��:=���� ��M�R��7�1����CQ����w���wDd�vacc�׮����������H��e�f�T!	�Ŏ:r7ߗ�*����vZ|��v��uS�VTB'Oe+�Y���&��tj��W��E|(4�P�}��5%G�@�H�IPv<�l�H[�y����I��?�8������؀�(��G�3,Z�4�sH�"Lߌ���g�)�%�T)s�K��������N9"���^$O�K �ȩfd[�K��߿��� ��"M��+nH>"���d�J�֍4
����iʼ���^D"i~2�U��@䟡z��SXĨYU8�����$ѯ�^�֩��[������X��:�AIΨ��~ �r*݌�eWTT�)r(����jP��9Yֿ�sd��w��$���Կ������Ɋ��u�AN��o�N�|5�!�L���N_F�<� �^��N����-G�"�	Enpz��	���C�԰>�qҤg��s�x��8�����B��^C`˷O=��w��s�7sH)�'o"���cyd����>�o�=H�L��EL����@.���*Zt��u���
O��
D8i��R�8L�?�	�tG�2`Y��\!��̬l\77�0V�����` A�C�E۱�'5�ق��t�[k��ܧ��7���f��{��Z�2]�2��o.>�o�s��'���?�a`K�>�����'���LphhjV�U�Tci�׵2���i�R��R���!G[$W�9Ǜe�=
6q���A�J!�����uwf�m�S�,(�A	�� G��S��o���C-�����pqK�7T-�۱#ݰ�����1~�[:S��U/^��s[�R�1�8������/)���mh$t<������N�tiޞ�%���EH2ZoI�m����y3���N��s�	Z]iiiq��������<��Oojn~��6۫2ƞ	^S%$"r�d�����<�z)��e0�f݋l�]])��$hJ0a��S~]�377Ϲ��9��"{u`:ߔ����k�5D�]s��0�c��\��ʘ�ٞ�bG���U���G��+���G7v&F/v�X�MKK�`V�=x4x_Y�W�5)iim�L����":C����ONN�1)Kc�,3���
��F�[iG�A��I�����G#�,�,��֠�Yg�}XChO�ϒ��ӗ ︈=�� b��lM�r��_���9���t-e(hij��;�Y6�G�!��|@G�^*ڷ��pk�)�-�m�p�X�gM�y0|T^z�.���A�%256]�L� t�W��a��?*=c;�����r}G�j\�g���h�:����$\���=�r �>�;��'Mvp�s�=���ZʿϚHm�MxjJ�F�\净h�#�
���G�p/�d2�����K�M[swRt��#�#���{�����Uu�����'�cU�����"�٬�Ax;ԓgϲ�TB�)S������a['	�;Dwt�� �����\��!
��w�|'�9��ğcO�<��M��V��M����D���v�{>��qT����kdd{ҾW���#:�<�o�GY��ԻQ ��6���77�\�c��SJ;D��鮀X�|��_�͐#�m l"��`EjA��N1�� ������Z��KH�R(��kK'r���1 8������:&���3�7�Ϩɋ��{���/I��M�=(_(f��Q9�4�`P�BÖ͛짺�!�UC;*�!�O���y> ���r�2�9�V��?����I[�PX��R�-TC��g��~�}f)G��5]G��M�ˎ-�]��hD==�D�����\��;v{��{����#<��FGG!U�͎S����m�hE���D���l����]V����

����B�`�[*�HW�}��FG�5�?7�4B3s�pﻏ�$�&A�j��1$ X1h�I��Wƶ�4t���6���wM�ͻ�mll(%6d�� ���ޣ{��V P��w���5��!�S?�~���}G���|�ʯ�DG�X�p����>��V��T<
��Hz��@�z��{�DuPׅ�HQ�g��V >}�A�&�)"���O��v�u��n@ �o7Ĝ��_���病L��Y��(*h�T�l����e�8��>J�ڥWXX�M����0��#i�+�:�]�ܖ����Ϡ��a�=�KB�ya �>v�^Q��?{��ǫJ�����d9%]y�	(���kZ1x�r����Ҍ5�ڔ�}��ȡ���@T1��ީ��S�p�4;o�ˊ���΃���o��oim�PU���┚�j̗/�d��X�F�Y��r�lm�{�Z�(/�X=i��ۻ[�A���(Ǚ��Qnn�فJ�۰6c<��g �7���,����clr���j+v���B�u+PhۉϢ؅{��cU?�(!���y�h>\;9${��o�Φ�s�2%�ˊ�w�w�>?(Ҁ�������[P���/{�TB�V�0�m�����z\@�O#�iK�� ؃ ����h{�
[n�W7q���m�����H)ߪ�"�r���.�pǥ��n�
c�jH�� ��
��vj�\�p;�j\����V���z
�A��X�rƘ�w7���^za�/, �-���p��ՠbU䈡��*�*����sNY܎�)�D����=�0������4�ʘ�nf�,���D0�����
f�u�;���f������4�Z��|(����.��غ��|�&;Q��
rk�?�ϰ�j^�����k��k�@1�@z��Rg�I�fuA|I�O+��~ř���rwwTe�D�D)���4j}w�j��}
X��� �^6q@{�r���Y�+�>
�r;��c��NsˮL���{u�T��Fe�reaF����tEAa�B|� !�����M;� qT9~�X�Ef�;8j���n�[��]Q+$<��
3=,��zͬe���c��mËSݡZ+XU5�Zߨ�b�Hڵ��i�����j.[*���*�S�Z������H�Y�(Q���ƺPw9���m�Q	#Q����m�iέ�7}��_R��,��W�/��GD+o��1i��j��?�igc��Ԅ��k�蠱�1�/caA�� >�D^�>��a���D���� b@XX�[��5�`��rYY����3�Ǘ/_��-����n��'�!("�.�kV�PГ�<)�n��r���{��Hp�h4D�J\�����k�Q�Q�	����f����>�+E}�y ���|~	�S���Fg��JF���Ty��k���y�Zv��P�lN�u�k��]��ʑ)�����pr�ٷkLv�������f�HI	o�`�a�/��D�|ن�݁�==�����t7?>��D�"(������eу��j��F��@bd^��]���$���Yd�_��͏����� �ؑ"��ݮ[�hmOR� �>à�c3�$eJ9=�Y�W쐋%��Ah}2"��C��N��;�恺V�Z>�C�N*	P ͼKY_E	X��g�m���M�W�e�ũ��n�CbU�l������A1JAˎ4�g�>-r��3����ٿ�l:�w��y�3���P�ǚr����{��I�[�?��щ����EC���?o$�N��70�Dz��m��ވ����Z���P�̝��9�x�����ꉊ͏wsR�U��Q0D����$<�."�c���S��&�-?;��߀�k��l��2���V��65��*�8��־�6��|������ ���VhK�9}�		����5ee�=Ӏj�/�{�f8 �X NmI?{�[)��EC�d�zy��%�B��?T&/�Vg�P���q6���S��߷���49e�q��<��:]Hb��5Xس������m�>O�p:(�Z`�a������hC�m����!v���h�|z~_
L+Ruŀ]�쉧"����:�"��O�2M7��".�bi�u�O/)9ch��Q0���=�_6?g��>�L4A;h��ϟ�Y.�?,,�!�6�����ߚ�I*�/�ɊQ$%=ۯ��Q�`�$�|||j���o>�v����u���yd�:�tZd٥�b���p�X�̅@>� �4֒���'���D���m��\~R�h��P*Z�DFT����=i���CM��� ����ێ����H-oO��p����ӢO�P�������w���1�h��KcM��q�H����b�9p�ya<����;��3U'�rO��X��E��\i�k0���DWn*:�&�@�&����i钿��`+�b#"�ȼ����W��2�� ��N����b��r�����^g���h�i��y�wšx�s�Ac���h����-������w ���e�s���D�Eԑ���<����u[+u���Qԗ����&ܤ��*�nk��Т��s�LN�f�&�a�S� ��&R�������{��A���h]�?��S���^��G��c�~�H����PGƁ���b�]�,�k�D��;vɐ��1������p
`��\h��K��3��l��{�����y�f>�qA���v]�b��k��"t� ��z"�T��`���<��;,��8�ס6`��N�s�U��KhFt�
�eτA��@*�^ȲK��R ]��Q�I�{o����������aIDj�1AA��O~h�2פ��,J�����̔;y2��ŀֻ��r!��'8�D�jy��?3�s��Ƿ��m}�G˿{���`����v̹�.��5 x�e_�6Z�ۣ;��ۖ�" ����P-�����*�Νz�18�� �ܜSRCdǽ��h�l�!���}AM�c_�5�q�"��dѦ��Y=gi���,q�c`UȻ.'6SCp����f���!3GF��U�P�;�f�W�}	�r����ય�xR�\8�6ɀ��o|I�_�`~��d��(��_vs+��w0���
o���v���X�ࣃA/^��:L=���2]o�kh�9��9��� �Љ^����h;ȣG4�su�;�9�@���+���,Y�4�g���@�*A��Į]���l� �J^B�5������n�� h[-�{?�?-x��ʀ7cjQ#GD��7��Q#M�\�*�Ch!
��A�����b�Xs6ZQ����\o��_^������_QFؼ��Q���Hq����A�5?���!z*��Zh!�1I��ǀF9Ks��
�2���e��]��� ,�_?�W�*�X9����sOQ3���n�͎V��@�uT?Rk���
_A}��U�霱��55�Q�)D���+�k��s88$$�ǣ�ƗM��E�G �<`�t��4�9��-��.��g���;_���Q ��4��L����.w��R�m�;q��Nl��X�doq>��tP)t ���ڌ��W�^M������j`�������,MS�BY�F�:H�-����T5BɐV��Q���g�^ii�?V1�7(	z���a�m���p�f}%N��I�0���e��מ�Χ�dh�{v�Cp��{��達�%���^6]	!x�vۧ���t��&z/@���f"Z��l?4t��՞��;�"4D��
G�N
�Vkg���@�2���:c]���N�m%�x�*�Y-��X#%�]�ݽ�֒����ъCC�w(�h�ҥ�sc�֧��p�ЮǺϟ�7�;N�k��u�o�Uvr�����G�߰T��$6����	��V����X����o9�ʹγ���f��d���t���.y�:�8j���|������oL��.��gS{�-Lt>��}�r���7�,��G�nZY��4kMT�~�ۯ��{��m>�Uz�??�T2�A����8�_
(fe$PETW���a*��Z�,�HF�-�Ϙ454��#^�/ٍ��=Xlǀ�ow�c��E��v<����4��J��2��d��N��:ZCAQv��ȉ�?��B=Rs�k-:thD�	h;������X��J�U��P�F���B��2):��٪ZP\�����x#B��6D�(�GU'��{�����y�'".C�������8���+�7j~>�+u��~���?�����a˞�f�T6�nV����D�~�좙�[�}����^n�&���� �Hu&�S�	S��k�?��X��Vp�E��96x:��fXa\����VP�Kê�4��2���	 Dpx���tcSR���0a��b�(1$(���~,��i5�zG����7���[�Q��2_�|���}U�τ�cc�(L�jev$*��_T1`��
(�+D{TE�"䂆�.N���8A�cz�*�	� C��w�Ƿe7J�����i�}�=���;�k<he����-��oվ�H��Fya��Ĝ�Fʄ�(ǣRIy����Jg�����s�IF.�=��I#�k��f�9�=Oƣח�544 n +��K�թ|-8g��<K�t�鞷 N��1��L�֣p�ͮ�"�[��H�cz����Vph�:V罡/Z�RW7ĥ��^s[��](R�u+y;@w��7�,��;��3M���������"�t�������={�F����;y۾��_S������I�we� )Z���� Zdnj��h�)��=����ũn��۷w4��F}�'�����[}����]#�	̞�:(@�X�Uh[1Z��A�I��P���~�rMS3���F9��عeW�zL�//�s��@^���~\��_�|��Uc�D �h�)��0� 2��e�8��I����<������#�Om�n�d�
��������v<x,s�����������/o�>��ֆ>��N��]���%��!p�˃�����4 �8}���U�P�V��HE狡�9��IQ�*��l��� S�,ӳ>�eB���=c�}tX��b�� �
����"���O��%�CbK/���"�/���rsHV�&.M���鰈�=44�b�wɼ��s�<�	�#�Ǐ())�Ra��A�M`����=zc	�ߨ**ꂏ��+i��^CE[<j6~�eTr2��aCp�e��]�����E�  ��l�Jt�rJzz.��"m�¯	"	r����֭ ��x{�Z:��Yw��<H)"��y���U�g�Ë�k8�)e4����N9�wpԤ'z?��C�?�kٽE9���9���o ��o��8��~	D�.����n�F��7�u�����,L����,��Y3�����׮�>�V�R��*'&rcE,�~�.O-"��r�92&gdP��73*��V@&8jf�S�}�'����7
�36�����x#
���uki�}eӞ^`2�v�ka]}��
�P+��Rđ��홰[P���eR��0���ϵ��"���|Ǐ�fէ��
Sﮮ'u �ww���!l��4�/ HE�l(7@t] I���� c���ގ��q^4�7��Am�X�һ����v����.�NV�#��.N��L���\��> ���i:��X�'��ο;�,0�����_a���ZUt ���7�`�o�v�l�򂉲��a���-��	O۷o�����	��<�^su���K?��T$��V7z�w�{ 8���>.���V���w�#�<80���}���1��5�|v0�CZBYZ F�j��IC{�x�#���e�ApQ�s����]t[1�ڥ��`8��� }��q߀:1��Z�x3�����y�k�����`9o��!x���$Y�����B�k���i�d��9�G�f�w���0�N�s��8�p�z�����:G�����//�	@"�h�:�Eu�3���G�^�gHQ�PS��q����ɼ���� ����k��5���������%���Xu���RnYOZ//-��-��!�7��G�����V��m��Ra��<O^�=ّ`|L��������VE'\N�����>����2�u��yt�n�nU��a��U�[���˖��U���^'�%��=ݶn�$��H�2���]���r_�8c��Ih�JKCH,�m� �Sw�J�P�q�ut�x_�^�6)*ly��qs�p|,�"������شF�9UYG���5�������ם1&�i���g���b%�,0խ�(�\��u$fA�L�s����Q&��<�Zv��#XXx%|���5�64)(�lG��Rߪ"���	��<n��y�{F��,���Y�:/�#���G}mՋ�Ė����I�%��9;;_i�Ph�۬7�H��U��ϗ'��U���N(��+���G���L�[��7��:�����#����{5�G8k���W�#w)����\X\4��)#�eor��틟H�+pd!Q�֣F��3����N�C���Fx�j_r��L�VNk`��R�l�Ѻ��e���b�Z���I�<+��#�ra�?�����V(c%����;Ez^��BNw�i�kY5`аt@�Rbw��#��g��Y��{m�10� +k]~�b:�/���W���%S��|���E���m�p��k+�)fJbm��p���uo�S�z�ﺂ�� ���4K�v$V�K�;Uw�g��hmm=!�;u��'��%�� ��!Q2=�w�*��?��I:�wu��I��B[���y ��˅3e��������k���f���9���� �yR��ۆZ��+*He=Yq�� �m翊�@dJ �r�s���}R2q��f�_?j|�tw�����kp@x3��a�+⧤EG�Ϗ�%m�\
�?^���9�~��o��/�Y뾒��"l�'�0�]��H�(���1qU�-�m��Tƾj<�i��'6S2�u���/Q���)R�o�l```U���o���6i"Я��vG@U����@hTT�	��
��J***b��?�;(2F����W��p��Tm^��:i��3V��I�������E��b�k��ϔ�	?kyL�g�+����>)��8�a��ߍ�H���!A�$ ���쁋f��`T�tJ~n�+�U5l�����?��i��ì�
Y��P(4��L�<{�r|3�������!.F�J���#�K�zN�.}��h�4b����t�����6�R{T���:��T_tT��1kͺ�sH�P�Ul��ֶ�O����қv���qDNjEp��3��0!����A;���G���9���̺��}?��#�$���o��TT;�P/�%9�lP�H����� ��35��5��Ut����6�޷�A|�s�"�|���������������7���� �����.��j�i���7�U^t<&�`e�č^k�����I�7(�r-��t<o�4��ܧS�U�!<˙�}o�7��%�%*�p�-�o����l�HI��̡����x�8��@�:R�I���|�R�+Wm~��xM-����pa��'�� �N�j�f��TԹ+V
ۍ7���-�n9��eX�`����̥Ž��ٓ&���k����1�%N��{���؎}��\Q��{X����ښ 3�t�qdfF@�YC�幷\"�����ǕՒ�����W:M"Ĝ�,��l��@8��D��+FK�.�"嵘
�>u����Ic��w�����iZp-�su��%���Z..,�.�j>�������5��BA p:�����8-$�����ϟ��	��^���=Cxzz�30$6�EmXq(�XTR`�i�a8��������m{D<�X�)<'���@[� ��"��������>�@׼�p�X&;0��d-G�Z��n�	p="��z*]��"�]�4#���N�7n�Cb�X��x��h���)��n%NEqq\9���Y�]��g��U��%��$F�'�zߏ�UX�D!b�������|Kh�#�P�Tmu�/���?zǍɁ�a#7'״��#���S>������'9�h�����(�+��4��~���b�E.c-����8Ϳ��8!�����i�?ND�j<8�}��a���*g��(*\x�<��|e�����O�I݋|90r�������������l{��c�i�H��E�5\o\�7qXc<�	S�\Z\˷q�����;p��q��xs%�����]yk�|��z�GA[�� ��������]�4�W���)���G�s�B|my{�b������O�����Ls��W[8o�v�o�u����5'>���h`{���Q�]6�� �sC䟤��ʹ��&v�s����3�5�BW��88)C(6L�K� %��e�`/�h�ǀ�˧�:_��Z�Bx�|/W} }(�հ7!��7]���ʸd|�<�Nn�3�82��w2{���x<sړ�>�>��*���ύ����G�Bد�x�>ٸhx�K;���a{��q��aW�sz�<����r�t~W�Hך�c[؀� �(�,�����<*O?�6�Q��gǌ���Z�h<���M��%��m��Q������9:7%K�f�Ls\�6P7`d�E��o@�ic$>���-�p�*В�<��;�ʳ7u��I���J
�}9���#\Yzc�q+"�vԈK�o�xe���E�K��'�x��RD.��ǵl�}�q���e~㢞p���ړ	�v{*K)���b��P���8y�`-I!>9��ha��ce���O2�\�B��T�\�����o��R�m�Ŀ�� T�C���4��� _� �{�{��&W��i�\0n(]�Y>�_"Ng����gl���~/�Y����F>�W� �����H��%�Η�w���o\��й�-K+�(#��Ԯ����oYr� '�=w�>y��+ܹq���Cwg,������4N�[*K(����q�ah%���_��Cq��8�	/��G�7K���A���wj���,�:�Y��������Y���kʴ�z���}�j�s�=��r����O-2�����n���� +0V��R�hrP�F�ӍC��k��%V�����+0��7�l�(��������h`��� F���W���z�ԇ�G��ȶ�ȋؼ=~	�ʗ�9o�Q!�lĽ��K*�����}�)��2�qEcڦ5�W��|��
#�?����%���vz���r�IxM�%��K�ϸ�������)ޠs��iC���[[��78��ytYqb���@�eX^�d^c�{�7�C��B@j (Y�<�Ey������{_߹���"��EW�Z�@6>���z(��8�Jv��m��k5��*6�n(H)�&��] G^u�ʝ?(�, �ٔ [�p2%�LǙV`�˙FW�����MTm�s��R�����,�6�xNd��Ӹ�G<��*7��!c^�Ob0���B0;�Pcz~ޞD�%������[�y{����ɩ?���궹����Sh%�c>�*R�����6�WU�T���c�
0�/�u\${`\�ڷ�_�f/
����������/Yg���(g������Eeٌ7��PK   DU�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   DU�Xx��{  v  /   images/378c5108-814f-4376-af43-2b942ce8b9a0.pngv��PNG

   IHDR   d   p   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��y����,�)��
,(�܊Z �GI,	�hJ�e0U�L%1��M�	J�R�T�3�VPP9���h)�*�},�f>��6������μ������ݷ�f��ۿ�����!fΜ)[6o��G�2��~NY1n�x��?���8?+D�;?��\��)��#�zFJHII���R�	I��$�r�m��/G��nݺU;v���]�x�ĉ?=򈴽�B5jTIEE��%��v�r���E^�|i��6b����s�*--�Ӽy�mNc˫����ֺu�Z/Y����W�Ąݻw��5k�w��c_��u�:�<b����c;�>iR�6�r>��1x8�r �E�i�9N��#%S�N=��<�F.���T62�a��'�<�Q��NYQ��3��9�f����(!�1�)��EZlU�R��^����A�WG5�J2�Ia��SJ%){2��Fd��ی��p@�*)��d�T*��#ED�R��E�MH3�$��Q(�׋��<�*B �ze�v�&M���ϗSO=Ujժ%>���+//���N���k�Ie�C�`�삐N�+YȨ_��<Xz��!M�65d��9"�7o�_|QV�^�uYO��N7C�R��y]٢E�����Bg&{��a9z���?��ʘ1c�^�9s�x]��Z
!�dԩSG��^iӦ�:tH���:�b�"{��e˖y]�9���k�����]���)��R�7����ǳ�̓���٫�J������c���<	)--�����SEQ�ڵkˏ?�(_~��l߾�Ѽys9����3�4�8و�v�ܹS���+ٶm��f͚�v�u�Y�$�~���ݺu36����~��r�i�����%�B{��5:���_��V�?���.��C��9�c�� �}��Y�d��\���q�N�L�/��cs3A�k���^�hذ��@&!|������[��
���V��-[��k��{�'�֭�ѣGK׮]]+�&�n���ɓ�K�t���H	Z0�PG���;��ݻ�0�|��9~*����4i�|���f����/7#�N	Q0��~�i7n�i��h����婧��M�6I�Ν��믗�-[��ٳ�wީv=��g��F��%�\�KC�"#�`�C�-��"eeeU��3�p���1c�L�8�|?��I��E4�@*n��&�:�ɲ�,����2*�nw�>ț:��o�p饗��9g�`���X��'�1i�'H*	������hmǘ{Վ
�9ʷݾ��/̍	��ǋ/��H�C��h���?6�$m��x�����ꫯ���7��Fʆ�>��b#	�*�+)��˗K۶m�}�" ]it��zm76���7�4^*��G@'���k_��u(�駟�nZ��i���L��aO C��\��Zto��v�Ֆ���7!0ML�Nu�,�B�R���Dp�>�CB�)3:�����k�8� ��i��@��o��+prpd��������?�5Z% �a�֑4-�7Б�O-a��6���3�Dـ������lL�.r�]wɳ�>��=8p���ӧFd���T���1~���Z�[��YP��~G�k�N�^��s�q��i�5�\#�]w�o5�{��ѕ�Y�f����FU�޽rH�I�'�\m&j��|nw�1��ЪU+әL\����@���v����܋������߿����&!
H��A��)~�^`�ѹ�D2��]�v�Ha��N��تhH����d"�\c`)�+1�1a���3�e�0�'�:b{x��5�D�Q�q�5.��l��/t,�'��v�Z��}��U-i�Y%N?� ��sUM����.3��IRν�t��t<���[I�v� �h�'7�ԑA���w׬Y#���Y�3U���t,|��}��f�դ���U2�>CCr� �Oa)����gf�I�g���L$bϭ�<���k&�v@G<���C%ԫW�HM�	�ù��Ő7n��x7\ADi!����D\���Q3�r�#��0 ��_~�J*�.w�ѹ�W^yŨ�+ې�O���{#A:[V��*�!H��J�B'a'�.]Ze�t� ���rIP;�3f۠�r�e��ұc��II���xhH���^î��� PG��`���
A�b!2P�O�St�ڝg��(��R5�1:�Ĥ2J��(	��ٌF��m$�>6)ԉ��z���G�N!��ݠ�u��E��&�ߩu>|x�7���] ܒ26)ԍ:~��r�W���!!�4v�1)������^@�w�J��9H�+
Jҁ���J��SG��Rg"�a���t��UU��C�6CUuָW!��`��0v��ґT��b�Pg�ΒCX��*!4�ap{��$U�	����ԝ�v!v^FN�E%{Αt(!ԙ����s��%�� .UWi D�u��ǰ���	A�"!^+|I�NbD�NRo��~�a%و���*!�%�����MB ��7%s�Nҡ6R�#��ik�Q��	�!��X?K���O��R�m��XmK�v�=M��z �6d;�"���:��4��(C�+*~O#������n��YZ숽�:۪���j{�¶9�����4�ޥBhK�UBX�� ͕�&B�)�L[R�RBpu���эuz�?,Bb�F�	��2)%	˶�@!D�m�-a�ؽ,����R��3��#ԑ��n�7m(
\�1�e���l�>� =⍄Pw�pR,Pi�&�鱓B�,����I�����A;�i��e	{q�E�MՐ�{�jr�:J��A�A���4�nCPUl��<���V��$IJT:4�p�����1vB����;��H��$0`�|��:S�B���e�H���yDrIA
�7�=n)A:PU�t�n���{oE��To�gϞ&�^���8s\��������}Xԕzr2[�h/#=�%I�b:��T�D�uPI�����*�#	���f�3w�������7����(<[q����cT�rE��Sn���;w�i4��� �&^�4jR�x�v>+ꂋK�	F��bY����� {��x:�3�l$���&���'�ãb��+��������DI���#�I��N����Lbt"��!�"��~��"dY-��h7ĺ�K�� 21?��9#R�0:È� ȗ�z�Ǆ{�+�zN�"�U2)!
$��4h��w��[�yMp��D��A�n^�ZեW��|�P��|�� [�WRDN��=4H�*��W^y�ɟN��?��H���O�#p��$�E t*���AA���zCق�6Hద�vC��a�T�#�F1�)�R�]o��B}�ad�&� �؉m�ӳ��MX���h�!�
���S�\we�����@r����DoI0L���u����r5ٲ�ѧj�{�d�9�[6<�6�m㶝MN]l�7d��d�!A��UMr�t���W瀙=i� ��s���g��7o�IG�[}�T��V��ɶs�w���g�0f���q_�|��7�(�2l�^K�A �#��:�Wg �*)A�҉x���r��,M��@a��R�o�Ѹ�^n{�B��O�n�`����$��_6�8.�<`�q���5x�K������Ʋ	Aru�]�I�sU˼�dj��e7��S�L1Qk��̭ ���ow��BCU�@׏9�*�;K���  Y\[�7�X���+s#�[>���g��B��,�# )6!
��իW/_���&D]�E�5b�Sݙ��v���۷ohG��阢 d��\^H(3y���O��D70��o$oG�#6�X�����$�n#��yo�t�2[k�	ڈ-�f!�G��(ؔ�7�z��/	��U^nB�I����T���xd�ʆ&�3u�����p��\��6}d#4b������Q{�lI��B�JuW09eՓ�N�lo� �i#4B�����L�e�'tm�n�<^}慼	�U&UA����:SwB9A�w3%"	��<+��"z��9n��L���zs�}��n¢o'�6m����f-=M;���6���۾�K_�g��C T�~�d���'�*���,��Q:ԝ60������В�k���|��T^���Z�bE֛R�M
��(
�!<v�X*q�H�`��Y�l�R�<	a���*[�� &��F�2yߙ�2�ѷ�� D{yӥ���$�������B��D�N&��jC*�wx%��lR�I�T���-S��x0�P�+t=�]����=m3�l� '@�8�$��
�(�:�~v��BV��-�0�Ÿ��F�t���ZM��o��m��L	��Z�m��K/U�h�p�p���4kxT،l�'�;(��|ڮ�4�w�jx�B�v�?��z4]IH/�hgM^�s��ľ�����g��>B�:���ד�����&��i9�'PM8<Lx/n��)SՆ���')/D����M�k��jFR��4�c�XT[�a�T��̎�-��L�l��`�S�f��������E��9�����?N��SfH��(����������p�L)�& �^��e'�:e�S�;%h@�H�z�lٲK�=���Ks��y۷o�$��,TtEYY��4hU�a���qp�ڵ���˙b]e�}�y"�E�����d��>ܥ���L������ɓ��r�*�D��Qr��ѝ��o+��k{�z�ߴk�v��<^j_D:*����ϙ�z>Ǚ0�csu�����M0ԑ ��_�����}��?aB�u���3f��M�r^�$�85�5�*D=�s���HH��?8`D,ȑ�    IEND�B`�PK   DU�XH�:9�\ u� /   images/5bcf48fd-3e7c-4271-817e-97f3eb0e00be.pngT{XT[�7����t���tw������]�tw�R�1tw� 1t7Cw}{�����y��G8s��k�������(-��N������A�,�4�ݑ���O,q�Q�_wm�}��>������X�)�"!�5#�Cn5��?$�V���4�sж�Grpp�3�0��նҧ��1L��!!=C��^P�1i{��N~��d7�A��W���	?�<�<�qziX>}|\b���#DC�(셟�����@\d�z��/3��v�?i��KD�"y?�@�
a��^0O�O���q�{v���/�[E�'+�UH�j[��Q�r�d��~�>t�ɺ�s`t]�,m	Ѕ����G�y�S��O���KG��J��!:j.�:JSg�ы>��P�<q����f�6��`9�|FM{3DpM�N�G!���|HT٬0'{����X��}���Y���ꗑ�C&(�^_��������]��O�4��3}j��'pQ�N^�=�Hz��'�`�E1��Eo��/�s����$Ovt��������-��/ɻ�^��A�P4~[ѯ}�`
����U�,�M�Z��A_Z�3Id[�]��M"�z�q�t�X����,B�y��s���䵆���N���ƺ���f���Rv�1�54aW?���ȁ�u����,����m��ej�ԎNs谰N�Ƭ6y7!=�[��oXk�(�Mw���۞�Tź74]7={6�.��s�<�J���8!�u:�Gɀ눴���߳&�0�����Ⓞ�%�/P�a�HRR�����!�f��ޛ����	MVZ�R�����a�A�M�#�]s[gJʑR��Dj���[�6��&�y,��n�e��p�$�Z�Oe���}3T>$<�W���XW}dH�FMk����Ɣ���%�}(��pȉ��u�&R�ߌpg>�Ki��%��_+y�4�
�FB����>v�psȩk$4J¤*�"��4m���MX ���UIj@��c��SO6����d��GS<��l��2�-�/>�כ>���Y�%�t|Rz�-� �p3iA�I������D�z=q�bn�T*��uY�t���I���=>u����Kص�`�v���LK�	���7m
Z/�綟����t�8����4����Pq��<����Eb��5�`4�I( ���_�~Yk���sSAQ�l�zb{b�����L9R-Z���9Y���q�8tyf����O�9�S	�%bR��̿������H���u�޽'��ﵴ����ppr.,.~)*�G��Ш���������D�������]^֋����|��F�K��|$�p0�nc��J������*�$�S�L�2������g@Qą���.��'.W���HF��Ϗ��˻��W�4L���Յ4q�������?�r��@*�4V��chݵ��~��O!;���	��L`5��H����.m���U����ł���V�趶�t�}�̆���T2)˿s��5�-��]>fTH	��qb���9���>��$g���<88gH�K��܂�X-N�wο~����D2S<�0�����Ô)����)��&��ɨ7�f,�b��}\����l@ݷ���I���f.>�%e<]����sQjܼўo�~��k٩�/��B��8������Й,3vtv�ۼ6�_��N���c�xxx�����5d޿��������7��#t�pD��zo^�u���n�G3(��]�-E	�7�lll���zz/T�A�}�ߜ�V;�K��Y�z���x��K>����r��ˏ�qd�ѯ/2��eC�'�R�|��N��9KA����]���C-d��xL�x�����hk{{���Ooo��D���ш��dy��TE�˩�yՕm������I�m� .IЦ9����PU*-���q����_�����Mu��/P�,���+Ҕ���+y�,�v��}�	�ڲ)���h�h���ݿ�xuue4��B�����MY]]�=�xkPd���VmӾ�����(�q�S�U��wh鋫�"`3�٢�d,��m�b�M�Kv5
T�{��a%�h�n�O�D&%'�󺰁A����ۈ���k�������.Ov6f��s:\U�1y|^�P�;�s�D�~`)��}L�����FG�G�(x(+P�'O�UZ̬àT35��ﾡ��-Qnt畈��_�N�u�{��Qe�D���'�zpxX�S1U�z^*��J��XY1�r٥)im�p<<<��*���fS���1%z�O�S��!/�I�] ��=\�mu���u. @�l�ܔY�	�&Am�$��ۤ���������@23w�X�h����@�q]���7jH&��G��4�o�/�����)5$������_ %k���j�ŀJ��:���6��$9 ���X�>�ȿ3U9�>��|qu0U<�N��;D,�1AH���9Ϗ�r�/Ҩ�̡��:Yii�.�6Z��o1
��򔔔���.u�&�f�T����≄�Ik�?�O�g���w|�rs�k�7�\f>�0�H*��Η�nip�k�興�7��|�_�Ǩ{/�˞���0�>�kf$��"�WV�oo���~���t�LoS�+)�E��0�4�-b���ˎ��xٸ��9�V���z&�Z+���Ue�[�H�8�����B��`}�ٗP���z��RѶ��.����^��d6s��WRLu�����b:N�����R(���'>>�F�"��٠�b���7h���v�׶���؏���^�=��hH���+ 3�����H��1���_x�__�^�B!ָ\ۙݫ��_"����M^�/��&���5��%qF�b��ED�@H\jD��s����LZy�!Wœ���o/�n%�s�x�V,��:�_��sn�P�A�|q�p8�F]�=,�	�`�L���c�(���/{�M> '�+, �	�n166v�9_�L`��#��(�z�ăH����w$�V?�KܡU)Ӛ�s"��j�ԑ�9��`2��:��_ZR�|����?1�{�z����'���GZ6Cj 	02�J�`3�(��3�x ۆ3%���a���Xq��j�t2����8��h���8`5���œv2 {������P�H���W~O555��Ԑ�NO;GG������+KmC�w&���SL$n���ou���i�9n_q��w�<�2��N�&�����f�G&%a
XXЍi����on��I߸u�Q�����z%���L�J(�ItH�a"i�˨X�Z�b�u#���J4xΧ�~Ӣz��U(����[�d��@|���0Y�u������@�|��������0}�BA"9�aC!��D����aj�z�����O��c�5��(m�E���Yj>�AI�NR��IӢ��)9Y���5�
p�������X�PF���o?�^����'�Jl�F��j�.�@e��Հv!�0W/I��u���:4��Ld�W:ZQ�	�M&�Mq))ʿ�}�;7腂�a5�ԟ��!�g��X��3rrrh�uf"�auQ1� 4ݏ����A���9�_@�ߖ�Ek$.�vW��o�FXLLG�7���?�(1qq&��ԃ�S*�2����J�<����@27!�;���'w���d��Za#�ݑ�{��\r��q�x�3�H�r��ݽ�I�7Uan6SM�q28���������ρ��~5�����0ˇ�ﳆ�:
"�O!�ā,3h��^�^K���z�ku;�Q�a�G����o�\�z�T�Bӯ��rp*��ͧ� ���ݑT݃���	�4x��cx�ED��Uʌ�m]�)`�� �[}�D{��qXB����:%j�J+�	��VY�κ���r�SPxc��Pa1�S�^����­࿿��]*����O��+g||}}a%*u����!+m�8���Ā%|DL��ȿ����.��V�S�.��c����3s搨���҉2�~�A����ONNN�j�MA� ���}���O���r��9�ӆ�, #}�>�t��R@Z� ����;��q5ސd�i�J�Ѐ:@�w��0qG���db�X_7r>�R�?佴�C 5u���3�� Bf�}~2e��9/��V��f�RqST�ǔavxrb�=QD�>�~=��\iA
*��7�x��������?���CB��<0}�����>2.����ݚ;h ��J'�,%�	�?B�qc1ɠy{��������۫{}qL�R��9O�z�����(6���w3,��J/��oX�~#;5ƿ�!c��r�rc$;�x���/��D����o[��,�%_�=�Qe������W�� ��Y���|�c�>�lhh8R
�����M$ྰ�DS��(jYZY��Po��|�i�OV�N�&�����P���2����s��2��8<Z���{?U�߂I�6y"���?lO���u9�[��1i��(|Ĭ߃+Ǽ����\@�T��NW��x&}��i��7[�
�S"�Y4ݎ�"����, ����^PG���Q�Ĵ�$M��>O��R}��Ӆ<J���q���}d	[4`8����g"�g<>�ݒ���5h��{��.Nw)By�9::����F��s<_��%a{C�+�ӂPO��}"`� 	ģe�����t$�8�S����§����2�fc�},�L�F�?�O|� BFȶ�<��-�e�!�	S�#��h^-�������)����,a7���<Beɤ U������]���	{~iIf��U�kDQ�M�����JȈ�=�Qw�X۠�*�٥D&0r��5���4�5Q�N�uU �IWK�@�d�u�׬��t�h9[�D}\@�3��y��D>�t��� H��`��\�o������� �P�s^����7���x�`�����P�-�]�x����Z[�1�pT�Κ��͋[C}��e�h

l��
LL� �?�8�m*�6fZ���䍚������3�u=H�釩�/����˗/��k^4�e"L�	J,�B�gjʅ�B��":�IH���]���P@�Az2خJ�ѩ�����^+�m�Ka��� ;;�=r�㙱�)�_�4�emo��?��Z��餷��G�hM�X�C��S��}I�{h�JEKXV&ypH�=������3칐���z�'DBH�UDђQ,ФH��2�4�����p���v������j���&&��t<�q�ջ8�矋NϨ�<Y�+���r��z��`^T+������B���I��9�-o�CM������E��=�tj�5�*�V �@�O���k��N��M��{�" i���"�8�kxJ��@3�@���Eɼ��ϟj�p�s:�J�ZՕ��6:�m(�-����M�i�wP\1�yo�������i�32� �T�7	���]�_l�}��Uu<v�>|X�7L�H�,Mi����v�L�c��F&F��Ƨ��b�ߔ�7��<Q���F�/�8k`d�(*"�4������K뇊ѳ�/o� FFڀ�l9�;ď�px����}\Vk
,
�	.�1�R`� A��6d�"4��p�|�B����΃�^B^�2�_��`p�гCO�w;�������?$}� ~J�(����Y%G��/���򏩨:w��
�<��p�C�Dw�5,�:V�N1W�H!T:�?�Jt���u|��������Q���e�Ar��Pt.g%`�RG�Ύ�vm�6\yG�PM�BsGE���-�=9�ZS������T���b=�n�ר�v!�U����j���2���,w�#*����>�ټ7��V��?�d
O�F�s<�����`r��*m�߲��|>�8�����
���Cd6�dy����0[T�B4�#W�~l��]\�{��2<^:Uj~����:\.�(,��6�)�����B�{Z[� ����؝����;�H��lX
D���&�@� z/������K�Sn�] ����Cw�O����U��	,���>ڿ�pjk���m_��î\�yа�W��3�T/�M-ZX�g�.}�ޗ�] ���322Rw�<�uk���}��fx��9�b�?�񰣽��n�P�Ċ��'B�����&Z6�f{߹�o�+)�j��r��|s�9������e?��q�E��������j7U���Zj�%r�@�~%���������P^�^Wm��Ӈz/>)}hs4O�k́�]\�T���n�iYm�H��}K�`���<z�V��x�Dl$����Z��!��\@��r� ybiiY���d(�ռ Pn������� �<���n��uZ̿�L[[d��VA�}rY��:Ŭ۩z�F�I,�ZR��Ǣ��&C�ϛo ��,5q�ſ�nX|CS�S�����SW�Ʃ�Tu9�^h��/��/A�;�0�А;9��ZFU�\�69B�pvg�\���Dcrtt;�U-�mlJ���hX~*C
���l��ULL{#�r۳A޾�S��@Lh���J��� %�x�.P�U�r��ttt��)���/��ZR�%���CHI�[�a�p�����͑�>��*��rt���(7�ZI�2?�(4{�4��nkOչ,L���K7���B�D�Hp�����E�����w_2 ��և�i�jo��|.)���|}�u@J���oݏ8��|d$�ġm���n�ި���~
���F��R:Z�@�SR��PQN�+�P�"�F>`�~�t����� f?�~��$^�^n�D���,ƈn>�&h6UѿM�G�"����tY[[�Lqm�,��Z�o��+WJs�1)3V�{l�wr�P��n�]oM5q�����؞� l�����;�o��f�JU
�O�ꎆ%�צŽ�󛴴R�9�3�X���L�|�4H=j����>[_;3�a��h�� [�E;�l������9�� j�7Wŗ���W/�����uk"��Ru�����ʟ��Z_1��<�߃h$�7e�x{�yE	�B����Rk���xQ*x���}ݎ m`�|Ǝ�%�L�ѩ�{�̫�sqC��:
�0��䲥8�
e|��J���9w��1o?C[Gv5��5����h=[��Mf�8�ӯ���������X{���K����r$���<
U��ޛO5+++�ۦl��bW�K�555��d�[�a圻�a�eȤ�pڴ�g��}�~�JD��0�����g\�E�g%�L?���f&�L�h˛�A����`��(��	Y #i���G�3��Q|��NS���2ᩖ�E�0X<B���_ڵL[�>��r�cY���CLzq}fT@����2�G�j��œ;Vވ�5�`�S����v`1���F����HRtclXT�)�)��R�j��CHD��x�X9�.���G#��3�]|7g�����|�A��9|:˿�<��K,�FY��i�7�ް��1��LG7P֐I�[S�2��uW�Q�Uj���f�+&��%d�P��h�[� 𮺽���hi��F*@����r����j���s���g3OP7pT�sG���@|b�������R�6.�uu,�3�22K�]x�,'ˣ�LNv�R��e="!1���X-�$[��1�UDIa�=��o��d��z��/�����:�0�֗̍���d��������tD(������g�]�;(�T�)w����S"6���Z8b�D�Hc&̹1:6�s�W�9 &SGsn%�fG�%�"VO
�_c���pK��-KӮ����`���O
�̆���]��7�q�B��ˋ��S����&U5����o����7�
�u��E}au��"^�6�)����3O��J<�A&����&�<j}��{��,,,�Y1?��:�l�Ӕ@5]x�ݎ��o��"�';S�O	�%k)�����F�B�yC����UX��]�ޢ*�_����MT,]����� 4�RianT����Ͻ[��4���{�]|/ﰷ��sߐ����R�AH"�����63���; FCτ��Ҝ�<�dNL�.'�M�Nj�Ob �M��vl�*���u�P���3�j����J�౳�� ������z}�9T�oS:����� w�wֿ�"��d�m�����p��������5b-�CK�F���4+��5�>����g Ps��(Mл������+_��)���=�6���|�(���%T�}����q���*b���vg�5q�L�h!d���EGM���|��nEZV�ܴPe<�ܶk�DQ�[�Z-�O�������ҥhE��f�N�6����>�W"A�ame�sZH�*��ې%s�f|��Y��Ҏ`� ����w��%uu�7V]aR1����~}A�5UcO[Y����[�6��*&�u�͓T�
&x#ie�`:���l��z�k�A�Sf��✐�ZjP����v�P�jk
�h��bH�����+X�,����J�tľ�w~��YhK|c�8p�u
.�׼�G��A>`�| ���IBvf�H|M�p@7CY�$��tv[�3��pgQ��۞�n��S�r������Z�x&TMMM�����־���4��8��>�n}q}���ݖ��R�0o:H$���7nXPɤ�@�QUX�$n]^<�c?	� =(g���j��-яRX�V��zJ����6L�>�AR���0���jj��l�p�����]���Zڶ���@�h.��&>���)�W�kl_�\c��
Y�ث��wx�h��;G�w��6	x;������B�Z��T�-"��{����+b�i�(K}�M~�l>�󐹾8�*��������n��6��H����';��k�헣s���{s��=�C����
�_��(!ad��;��W��<Ez��-�[� S2Ay�a��Z��Cvg���F1�� �̮�E�7 �K&XM�&(f6�f���;�0ac��H���C:QRc��6#3� ;88����W1G�ѓ*����f�/lN���Yo +lA#��#r��᠞�J!���/��v���w��������G_�YXT��l�lPQ�"�v���Qr������0����QI'1�gE���"w?�c�F� �W��3 1˽9V`��?=����t�y�@g���������9^R��7��
gڧ��Վ�����G
p��ɉ0fg}/*j����Մ��������Y�=j�G����!�`bvDc��$���K��e��\�θ��l ڥCS�����'Qv�у�Mͭ��LLJ��9:J�@;��.�6��Ɲ��R�3��<V� u��-��õ����3���"X ��+)�i����4�_�*Zb��}�;r�}̡��t�����J�Jtƍ`���x�?D��|Vj�_�r��"�e� K��x��s��k8��P�N�ɨHE�GD
  F�@�ON^_�\	�ë�hS�:v�b�{{G�+
��PzRtD&'�.q�r8ȟ�^�÷j��f�"�DcbĤ�]ex�q�k��}f�h�:hK�oB��3[�@�gt���fe-5��d��70���O�*�<.���)KA��I���f�x�liU�� �,�������322dG����6�3�qO[f�c7=&��M7�5�,�.��Dt'u����8�Yy4N�+��>ފw�h?��Ksd�����g5�蓦���C�3�Ԝ+[@�wh�B�Fpvv6�Ӷ	�M�����_���� w��חX���-F��^x��}��ıUr�-��[2��X`P�'�+k{�����Z�	u�jǇ���T���嬢�jr�މ����G�����}�9�($�	����5\�S�b���^h�.,t�y%o̤cL�ы(힙�f�ݒ{��ξ�`D�b�`%�D7��]&#�,�=j�D$%%K<�2�ω��'- �ED������V��u�P�t9��sD��Z�cxzt���{��A��j��=d���*lEF�H��$M׽PGt�Vz�!;D@ 1/�tyzz&�a�:t�*{�5ed"��U�ke��(��0/�|�%̙�b��T/$l�pIӀ%�Ҝ|*0yD�0�p�-���W��J���@gk�ì?�3��ݻwU�����w���L| �����w�'''bw,��?��7w�����*̱r=J�f�n���&����u��������,/=�h7m/����w���(��pu>n=I��ۙ���#`b��0�}ʟv��+��ߤ��U\�I��ё��dy���d��@=&GS+❫ �]�2�3��c���eh=_JYc�c�R[N���JKr��=��i[l8�"�1W���V�b����f,�lq�#�Pw]���>A)�o�ӣ��q����A\w1����A9���L�P�M�Ԣ��N��v��>J^�Ttx�gg�l�]��Ӻ]aa�^PP ��.I9*��j�iZ�И"�?���2�All^�R�s� ��Δ �(W�~V_���������A�"��;I��д���~C�Z
���/_0��L�h�<���L�u����=��KL� �V�~]���:,� �1L��,XR�$ 0 j���иFJ�ԅJ�H�����M?��8�hY(띐V� %��PH��W�����u�O,�=]�j��ؘq�[�%JΚ1�1���;�����q� ���*q���g/'R�۟��sf?�aL.����^������a�R(�����6� ��bQf	***�{M�d������WT�<�A���4$����:X�a=8Y�w�k,�ፖ����,��,�����-�����G�8����
���I�m�XU�w�9O�K�����4��]݁�~V��G��K�"����m��_hNU|FIq��su�g*'��0'��|�-0�oc��$H�o�O��A��%��gK���I%C�X;����/�GK�g��@4τ��خb&s�/}n�P�T	"�&O���J���6WeI��]{`�Sn:�T�� �C�4�>}z��e��8]�)a>e1!��,F���T�j·�ے�d�g'S��nN���~!!�-�0�k��[<]~�O����;T*(6;��)��U)3mmiQ�� ���@�fjS��?9<��$0�M���& �a�G _ v&�M�8C���#���w��l��0�!SW��\�,Po-j������DSC���B���Z:�JüP��B�9m��!�����{1��yN��f�u���S�LdV���\�qqJ[�3jNW,�����/�K\vWi�$��5��&f�� �����0�� ��П��g�������&k;�gk�D�D7��l�\�W�s�.��
5U��7e�M�B��ڧ*��z�p}lV��g�Ȭ����%���hf1�(��=¤���lN�⑇��R����'-�!t4�M��<�T�,E�6W��7ܶ��µ͊���l����D�f���Ek!;b2��u���?>��
����,B���?l�������Z��]C�>�S����z�}%�~S��$���5���ꈭ�,�D���b�l��@�������
p
�j5�����G={�fR���Y��|G(a�L@N��>w���G���Fs>�Oّ�����^oK�n<��z�M�61�)k3c�f4&����t�W��6p�>,SEj��6+�]�ʾ̅�e�~Ng��	}!�,J=C,��O`��v(L?�T�2�j�wq���}L׷�IӢ_�؉[j��J�~�>{W�w�M&	�)4>ut�'�Ux3�L(J��Zi�3]@�a�,]4��:$*X��f;�骧�p*��;�ބ���i�NR>�*���Xz������Dʵ���x���fQdnт��r�����Oe(f�"���3�N�<Dֆhd�.-Z$Q&GZR2C��a[g'�F���;'#�i3�6#BB���%K@v6ᅦ#YX �[��+�� k�J���J�붲��2���9��]���,�9��?�������--�LY}��­��hI�u	�S�l"�ELn��8��8L�yu�B�gS(6�j>�E�6���ݝ�#�q�6�8�����,�[Xk�N�(�rq�u���:9m6�ӳ������L�z�A-�Kzz�R'l�������p�&O��U���9[{{�W�|r?�����̙�~9���?�Z }Cq5,%2R�������)u��k18���3�j+p,%80p	<�u����5�'���~�wINHs.� ��nU$����wU��Bmפ�	��>��`�a{ U��A<+��^��&��'G�SPQSq�����S���w�,�������UWqpss*��+��`��������љ������ht8zkǑOI.������^�d�T:]s�`���C�B�f�	��RS�r�ޟ�;U/-."�h�s����
`|�S"֟8�s���y�[�T �P�S��h�Xh��XXX���tV����p��rss;�(P�*R�+��[b;(b�Ȱ+R;<cg%�U,�/4Z{����4���.'���.O���;6��!��)h���,Sȯ���l�����5^�@�c�&1]2j�Iq���KK#����9b�ھhY�'G�:^��L�ny�2#�?)d���};'.Ǯ�v1�AV~M}�prdg��J��V�yf0Ԁ�v�B�٠a�'y����֛����8�Hٷ5$���@��j�(�T( ���oG���n=n��.#��7s��=^2SsSqr�؈(��O'ե����p�\_�b�A>�n�_ٵ�QܢR��0����u���z��Q��d������`��7��P?<��O��^���[�\����q���b �$�lS"n�	��VքQ��p��"�W�3q2|�_���n$�h�^���
@��Q��S�jɊ��	�,��B��']Z��x!9��v�'GF�j9�X�瞠Cj<vTC�__	�~V�p�{�baAt�0_l��/��m(�3s��82�V�1�%x���{�
����<���ƫ	x�{�����P��Gc'�z3]b���)��#��eu����)Ns'r�ƫ����|�'g:;��>�i�e����k�>}���q&^��e��B$��x��ʵ��s:�a)G���%�U���ίG�H�^
���z�V �C����R�Q���X����3!o~a�ʩ�D�f�z<DS�W�L��t��_s����]|�����k��ֆ��/צU5\�S�8L�P��F	�����<<<g7����R���Qx�*a��ˑ2�@��@bUU� 5E��!��c0d-�..J-���K6�K��)i?(vt7��b- �2�|��TT�����r�Ƅ�w��]�T�:���VS�{�ۨ�e:N~pr�M�D�$H��c=õ���9���o�4��z}�<O�4��!Ġ?��8���@�[�R��Q7�璷i�S�����hwn.��d��"a�U���ֱ*�Ѳ�M�r,�e��,=�ޖv��r\rN�j���S�$���_a=7;�n<�3CGG4����4Wkbb�L���(Z��=� z��t<�T��V�խlm��*PB�0���Խ̶711	�M����Çj�6ߨ���#�$�:� ��p���&EM7����p�a,��l�UvO���[;i޷{L�9.�'o=�2�2g��kQ�r�&�E���jq�2h�[���?cڿ���4�ʵw�c(?�VL� ����� �\��"��S�ER��c8Jz���p�&���{Lz����EDD��LU����
��5����ޙ�r���[�0DDK��^�_7�����z%7o�k|ˋ�o�����=�`HfF����KuZWﳊ)������~��渿�������<��ꉌ0�DO��@uJ�/69����bᄡ���j���M0�Y4*^��M�5-$M��L)V��~�I�#��;����W��f*�,�z�76O\�w/�w]ꪝ�5i? j���`l��E�H�Qͬ��c|z*��P��[
<<f�����L�$�&���	�zYj����5�R��D/�V���\�(��W�W�.��R��$�ߢ�*,���U8=7\7��N���܀�E�̎
��حۨ�t�K���������e߆ɲ��)!�F^�?[ĉcR@^Y/u ���Q�:���r3�Fn����_�Fl����#K������-�o�?���zyyq�CBb&�N!�DŻƹ��`�ę&��c�X�;��CUN]��N&�����76W�o�Vn��Fq�z?h��(6���k�b�=:\�4F�lim�t�'I�c�FC�� �Y9�[��7FSA)cu:�0%�Ԋͯw���{cb"�n�P0�T�>w�QP~�ړ��������2h����x��Ȗ\4��#+��B2>�l~q��E���A��(Bq/��p���"����w���c S��� =����"D+�d=��a�}������_P1���
�����^\��\���/0�	�c��݀>��v�锌;[y=�3o�@1��t�twpq���h%�Ii�%w���^8�%�����;U/��]͋%��Ƃ�����s���to���mr�j���Bs�1��eO��J⫹m	�<���A��;�Q�P8	ɝ��N5<ӭ��F>�y�47>��sRj;�ؠ_SH��|vv��_}}�]��F�+-f�5V�>{ۆ#���s�/���&�!��uy�;�揳�o�ߎ$%�?$?L�B���\����H�:73��p��֞��2ә�,{RX��>�؈��܋��rp�b���Zs���º�-ࡩ	=��A�a<�\Y^�/�-��v��'�,�u�5
��o8�Z�K'��5=O+<�}��Qr��j�D����6��$ܐ�����5�;#�mVRe��LjE���%}�vضȟj������W�.��xw.��k%�,�����dyo�&�R� <\8~��<U+y��--m0��*��@���\R��i���?/6��=1���Hق1�{z~H%����Z���4<k�	W�jH�l�?�+ṣ0`OX��׋~F�=S����
s��޹�o�����+���i��0����u#"1�EgC�Hy��ڟ�`Q8�U� Nvdp���YN�
ƛUPQj�\�w�+n��c^Y]�b�6�OBF�9�;��`*`�>���q=(�҇{"F*���~���t�k�4\w���q����?yw���x��#�$f�ďm�tX����#YFC�����b�?[�������l�1-�&}�uJN��4���V��j.�f�=�F�N3��f%y�Y��Sl.f���1�)���t���XK�*���]��R�>_�Z"�-�������=t��7$I[��M.�ϘLI�\<ȥ���P�0I��"xz������0E��_�y������q
��c��X�Zg
����V�?0�}�R�y�J��x��a��6����I�p0��@����	�(C����l��_�ύ���/G>_9C���C���zUn>S�Z��,ś�K��X���mF)?=�96v�Nц�b����I��0��wD�����9�K�m ��+;�!u�@G�.+���=b�+�'L�9��lV+P�U�%��:��1֩�W���%����';Pc�#����_Y[�ck8[ E���|��t����"�v��M��[F�px���pM�c� �9���5G�Dl���,�2{)��������Ub�;��@H܎�G��M����7�AU
��C��\e�j66�Cqz��xo�@ ��"�KJJ� �(P���vz��H*�����+���r�/�&L�"�ĖN�.�I��t������'��.))���H:�b``@$%�8!#/�jm�`x�~|�f�ǭ{KKK@���+O+{�Z��'K�ZԠ��`�4�~�c9(/?*�c�P?��
C��`���F�J���z�ҭ�*0a�d����[�{͝oj��x��Ü�A�{x����Ԋ\v?�L+̧N�S�YC蘱ǵ���>l��|DDt���rb���'�~m0U����6i�99(���|�7�
U��.�_�Y0�����{G��p���N	�5���9ʙФ�����^�5�wZ��|��U�h St�m �z�9�`�'�Zը,�:�(xn��ѣ���%�\F�\6�Y���Ӻt�`b�ہ�����n~���8�>��7;��Ꮔ$�7NoC�/1�6�.�n��k�}��#��ӧǂ��~z��z�@w���<�篗_&X�p�W*���ݨ?h�lWKoH�]������ŋv�AR�yvj��E�?��*\���w�Ǌ0�Ϛ� �K沲�M|�L>����)���������;$6:�95uෟU�1�_�@�9� %�Q�x;��+�����E��g�ϟ���]5��<}�
��SB*#Wl��tmZ�xe(,=<޾;�C냽!�s3Yn���n��(��������2��-�1\"3��t,?|-".��)�£���7�<�Ԣ����Rf,z5���|~���P]�v�:�aٙk�&k�%�IڳW�p��'���J5e�)%�k�����Έ��[�ݦ��u��_���������h�IT�f�%Ԕ���` ��Z�[|e�pa����Y|b�S��O>Y��!�.���P�%N�㤥��q�8>/N)6�x�+���6�K�a���c�J"Ҫ���b'����}\Ӄv�����/~�$$��ݬh�����Ԩ�_rq���)��'J����L�]o~�
I�w$l,RɨkD����y���j3S�s,�7�S.�k>Uq�<�r��Già'2rr8���T�����~���A�}\�O�?��J���7W��I�m���ྃ������751y�4�u�B��V�ԕb�+��R�y�>���5�����'����!��l����\���t�iW��$��&��1�/ݴ-u�{s�� !�q:�[���*��qE���.M,�?�<U#B1�r�	'��Ք��H��5�R-��>$mɔ�%(����?��8X��p�{��%�*��s;x���Qc�n�˩R�qnn��r7NEk����)�V9����so�\PP�؃}Gzl��D�Q��N�Er>�ռZ$3�X<d&�W���=��I�J�H~�s�r<�$#�Ž���߱�����震!���]�U��>��
>ϗH����@	ID�vw{�213�wpە7�kb�֑M-.����(�.[=�*�h�3�����5�����T	�'U�9[2z��`ˑ,,@�i�V�*\\��޷����I�d���ة�Z�������yq�2�sۙ�8�t����>�6gBB����/����э�rdl�o@ :�ӧߋ��V^�	�~����3&����'��h:˰��h�(HKI�����Hwwww7"�)��tJ7��-�zf��q]���s?3kf+(|��z��{�W�����P7��ݯ���E�;���Li��?D�c]%)�:A�im��S�7ev��
Ӳ5�G�kM���&�"=N9�-*JKi�ڽ^����477����;"��i�����3��gӝ���?����x,f�|"�W.o{(,,�@��͐����߫��4���W���d
���P�}L��~l����:��z(I�U&V0}~�111�>���>�ڪ
$^�tmmm
**A F�nO�mB{ӡ��0�e$9���O6��srr���vv�������W�������{��q��_OOOİ�<�b�������'�ڑO��ZZ����� ��\�LMMaaqA;�@A����� ����D˫�c=���SG<��˦��Tt+��<�N.��.��Q3߽����[�^QIK.���`�B�M��`���N������c�N8���wO�oZ
P�-��_��;�~�Xb��d|�R�-y���r���1�	���bR�4[�ZYYU���\K��]S(�ʢ &���"ڼ�����֨QX�3�Җ� ���H�U:�h���y�˺�������L�2\��sf��B=(I����/^�\�3�_�ކ���=761!nkK7<2��v]�YSO����6.!�sA%%)�%%o�h�������I�ml������{����£�H&2��3���qԐ�E���@���~�"jKǳ�������5�ǝ>���l3lKXUJ������P4��0t�Ԡ�$z�d{{{��H!���s����R̳���D���ͫy%5=͋k����G�<o���w�q���n+�ɺΎ�H�'6�r�bU{�z�ls��T!��U*��)&�'�=0w�r0ǌ��Xx��@�@7jlZ�%����/.������k���Ixg�z���v��ta����ђ��#]�6=�<���>������|&�o��Wnn..���;���� @�ݿ������6D�{~_Q1��X���P����GOl���`�k����hj������z�dz��#�C+q��9F���:KI�Y�z���O�O6JUM��w��k��r:� ��M���cbd��C��PU���w�`g�_��u_%5=��d,5����5�ۡ�]��|	�&!q���%$zj��i{pd�n>wƣ�Lչ�3.�x"�����#���1f�����\�^l�^��֥I�ܝ�Tp���w�ɟ�c�ոˍ�Ye�=>��dDV�G���:�U:��� �]��}~'� ��s���]�%�\ٸ?*�v�xwW<�fnZ�'��	��/�r�mt�B�:�F�.�~Enpp?5�Tg�w�䯂*�����I,��b^ܪ���GPP�v&r&~ӏ��Pcum-��.!CW��x���@���ps2��v�y�0�쬝�������GQQ��(<D�XA��5�j���F�y��Q3���EEp�����p�Wŀ� XB޶�*�������EL<t���⠧ǋ������&&���,~�-���̼� X��Z��i����!766l�4F���#<͗�{{/�,ku�m	)8ʧ����iP��86��Wo.|��۟̇WgW��DJ���"�հILr{f<�(ݖA����@:	�<����&�f�H��p�ɢ/EY�v�bߣ��Ʒv���w�B6"q�%��O�S,l��N/�~���J��.�A�$D��t��}C��㳕�SUYٗ'��v�ZKK��몬;Q��>0������uv���C!���^鴢SWW�b	TzptTDI	#!11<��=N��Ŏ�������&<�0�RR�E�91�8þt���z9SSJ�׋���aA�ۮ�[^�;����x ��'�vt�9���h�?Y�5�B�����ҿ��,"&���ny]O��'+/I[Cw3}�,��r�k�[a�ޞ�Ƨ��f����ܘ����/ߛ���m�?Ci���R�z���Qo�^��AMM��j{z&���l�e��Qٷ_W��B�eU�%�ґ�$����wq.�� e��k��nr�ߖj�-j��>�P���\�Ϡ^o��`���y5���$ݰI��!ȱ�N\�|�����c�:�(�jy�uVkv,!�g~��iM���!zA''f�z+��b>-�Z"����f�wj�Z�)��.q�������=x����%�1ZZڸ�̨?,x}� l�)���%��\&g��S�����aWW�|�7���Sf�a!ii$�����PRɦ=��}��F��hq��{�����a����Ѹ��Դ�H��g�	�O�
6@U�� Xx������vvfaU�x�}!A����tڹ��|�x*^#�%�����	��D���h�}�¨nγ�+�wm`Z:�nԢr<��Ry�c��;�<X��0�S	��/��9��_ppr2b�0L��+5(C/��ِ/���_��_u$���U�7&��ʕ�\�|ǮF�i��!|pNr�.��U|Z�J����A��.��t	�����>���Y�J��꒒W���c�����D�2�u8]�9��������j�V&��t�	�5===t�7��&k�,P�WHH=�
�m�!5��G�4�j��t���)���}��A�9w�gI@EQ1@��*�����0����:V�������^��7C����/���#�H~~~Qr��\B�����G(��e���o����VS������j�g[x$1�Rz�M�ŉ�V��hyl@���)k�G魳jtisj��o]l�})�g РD��e�z��C�8s7�ԯ{�VM��#C׀�%�^�l�G���x�~U�Nm� `��)��R�q�q���3�y�D��(f��.b���\c>A�oMȅA�3�l���͇OF>�������������_���nhH���c����7��a��#P�R9쉏���N]��D�I${����>��yg�J�rԪ�P޽{��Œ����q �q'��6�vǧ{��T�]����9�U���\VD88�&�#��ģ��Ǎv˟+�8�?���v��1����|�* �5���<4W8�9����q5�/6��>�U����	8��&�Ǌ�򍕾�ܖ�j+_�ś���$�Y�>�z������ɒ��Np�'t�ab$,jW�GU]�/5~�_텞��Y�0�1ZE�Q���⢼���U~R���G�$�h��&?����8��ǆ�]��=���~�0�+�77� �S��Ie�q� 2֍�pP�y
������x���������� hR���{B��yy	�CTljy�����OK"��� %�@�N��)!AA ��c�I�����Z\�>���O��҂�u���k'Vi���i+L�sxѮ�(Š�nQ��g��e��`�G7ggg�GN�]I))8�����%��+B�XW�H8��y[JJ"�=q���>�}�cA�NQ�E���:�d9�F0 l�H/Ws�ǰ<=�����H�U-A����7�g��̬i.o��|�a�̉M{��0� ���vZD��M��_��*|5����.ү���6"���U:��SQ��k�����n���uJ��t�U9���t9����N�`X7;]�\�ueUP\<ww&�%�˽|^����
w^��&^)�:����P�%�	F����F�����v;&H����h�P �:�~D8z�`����N=�NV�ǳ�9`��� Qh�c��5:��KRٷ����g�������iK��zNn��� ̒1t����ԭ?pG�`B�r�D��η��S<�,-i�����Z��	+��Y��������r0�r||�gV������ZـC#m���C����e��`*��Շ��߯��x���=3K�\<ܧ��#�%��3������<s�}���Dc�Sc�f������* 95���:�#�=�0Ĺk�c��W���v�>n%�����69UȤ��)�[��=rs�Ƃp	-��p�����g`"""zcf~نԿ/T��=p&����
��w�Ĝsױ|�f]"ի�o��F�}���=����tC�:=��4���`bՍ���q&�{�ѐʲ����֖H&n(�aK4�����XZ��[�A��-�M����õ�N�B
�����b����f-?�	����F��4s����^W��/���X\$�頀\��q�'�3h�$��*����`��Į��2&>>���r @ #/yxx�q?M� ��BC���-8��9mմ���>���*/,2�Ǿ�)d�o%tMtj	x��[�����5�T��>���yj��U<�6�9.9����.� ����]Eu�-��jѾs����d����2Z,�W��<�t6�����=�� ��"A�Ļ'uEf�sĈ��mN������S���|��}��ыkk�G���>�����ףcb���W�i7�j�~�z��{4�u����������Āy'+���J����t��cu�U�ojq�$1��3��2#��
�o�����`�!��5�c��]��H4����G�1X�ɿde� !E���̡y�����'�(˭?�t�#���f��eUS�J�xA�4O&={.�q{JJ���)��u��@����G�**A`v�Oue/�����>�_�333��*]�4JvI�c�  5&�E^7��*�_��7���d��{B�:K)�����f�TU�ws���it��klk�����u�i`m9���Қ���GA49�������{�N|�ڠV�8����✷X��$�E��Ȓ�����<�1w���`��(���i��Ś�n���ѿ�\Z�}�岾~>F4��#{��l^t�b�R{�"kc�� "���9J4x�u9q�AKk���������-��D�(i��JI��'a�.ܲss�jhzR���bss�CQ�Q����bw�ͥL^�ܵ��Պl�~yQ��CB��ftjcr[�]�0^�ӌahh]8��bhjJ���l4�c������H������&<�U)����"<P3�׫袨����8�^�U�+++���&�ǩ�PN�b�٬g�!abb@�*2�;33Sc��ܧ�����S����H���D�b�n�x���l�_�cUkM�����֖����2�Ke�\8��n-/&}���4~�1��yd�X����x9J>����x�@2jg8���D�%]�TI���9��67�}}{f�F-(�a���N�,��z�}�r�%l��w���*5����-7&++۷��ọ����aj4���w󨹯&յ���K�r�����x�^ׇx�ļ� VD�;�7o�y@�K�$DA�@A�	�>����q�O��������݉B�XOO�"ٌ��Vw�	 ��c��#M�� !�N�E)xOLCC���R�b7l�0]�j�7���1��<n"����g޷y�r�RU�6�RT�HKM5����U���f8�S/�D�d�'��\q��2:�b�t�}�?�]gc���K��.���¼�x�K:6//�8\diE�4���))_X���6�=5w��a�;�	Fn.�bI�iv��ݾ�d���Zɫ�k��6��f�t#��:�И5���i��U_�g���\p� ����1(9�UU�m�[-��	�����h�x%�H���=�8��Re^9jcc�h=��ŋk�3��f�F�yi��;�.����Y���Ұ��*�p�'�^V0�>g}8N1�F��L�"�cl���M��Q��1N�����7F.��R�g��}��� ��f��5�h4���I��@ʊ8�����y%E �Q���X�d�ے�/���d5�ߚ�t�.?�������qa`g��
W�o�����59?���B��P(�s��c�R
��#l/��K��a�7f���[�TT�DLŽ��XtT�O}��Y�c7�u7���%5l&_��@v$_�&FG'���:L��2�zw��>��rb�����:�v��+4�Íe$�X�����ͨ���� �|���Q��O"Q����
���p������!H\�E�.w����y]~���$$�"�!�r��v�.R�db;�'�[LH%�]�sJ��\�k����h�be*�ԟk1�|lX�lD,f�K���H���8���x�C�)?����6��x��v�����/z�O�m#|������DJ%�O�w|����b���EAe%�LU�q�k�X��	��BB����I,o� ��AB��v��'��1��c�����E�9�=��"��o�!  t��īB݃�E�����-�͙������X4`πh�3t���*�";�,y���.�TW�;.��Oױq�>Ř5:0sa��H}u gaa�F�ͤ2��8�t׷^���������5u޽�������_���QGŦ�������$g�5��ӱ��q���}����?c���(=�O��S����f���r��ϟ?���;0�>-o�׏�[5(8<�M��}Űں�o�:x�u��\T"L��f�$��?��pwi�,O�ʪ��A٧�8�$Q����bbb�����G��rMޑ�	mpծ4SǾ�3.���h�p}Q����a�����aA���n�i÷���nCI�/άK�X����2~�7��6��.�#���f����|$��ĳ���@����hJ�Xjv���%��������щ$���Y�gޜ,��[�� ��\.����m�5�7Y
)͖�[��'���>G��lqf��L�kk���@}�,�v[��f��CR��ܪ��޹TS��� XoT��A7¤�y�C�s��`B�Z��k �m�J��ccck49���+��%$���%�i��Ka���C���l�����kSSS��s>��迫����n��FQ�A���	&G:���T�ٝ�P	���9�Ɋ��> ]�����rZj!�F�jTr��kS���J��W�c~�/�/��R<�py(>&G������G�$
]�FQV��)����Y�KȖ�bO�n����g-���Ə���ɥϟ��-�ìm� �����ˬ�{��|�!��ul<���Ɓ߫e�g9�&Mq <����k\\����11��yq+�%�ؾL�;�	�d��B��C �SBR��Ǐ�D�&���ħ����)H����Kt��s�@W3��ZZZDL�Yc�FI�~�K��J{��Y���|��CTD�X,q��0��*�V8���mə�!y�Ri 6�M����L��I▱!)�o�lt�����]h������$٘�gcJKѷ;����uts	~���<�)�>pDp��+3z��b��5��Oʅ5sb��k9_>Vn[[-;%�9u�()b9�"��c~�S��-�����O�`Ĭ%�Z�z�1{(�R���,�7%�5i����NN����Op�A�F��~���ج�OM�yy3=*���	�����E6S�m�C��8)(�NF�����Y|)r)@A`[��DY	j"�mKg�@��,���9�ۡFI	��������!��٧.�f-a���r��Df����qD���\v�j	QSJsg>Xݣ��H�뤤$����3F�QbΦ"0��M�Ŗ���K��*�CFѠ�]�:�g�󚤝��#J���p�D��#�}c;�W�Y�j
�����L�"�%���ڈ�d����=�ܖ�i�ڕ��#���LLL�21��@���RPS#FT�����dz,`�/�Õ��	������Ȗ��,,��G�B	��΁�����0�}��튩�h���NY2�Y(y�GCԫ���G+<�D���4R�A� žXȘ��b�E�3����q[Gɏ�w�d�_�`o��A#����N>�ߩ���JKnv���E�#������N���=w|;Z�^{D��*�V�ؘl޲x�"�I;u)��c�"�me]�hP4�������|2e 912"������P�q;�TF�a?D0TU{�~��x~~��z0}.�y��"WII����Y�����o��'"2_]F&j>�5pk�,fQ���sƳx ��cr��eƍ����\5I~��J�G���9���qi_�mL����8����v�J-��lI�n@�B�h"9�)���`;bQՔ����p��q��bq
������-���7�q��<��	�&]Ŵ�4/L�5���kim<PO��nƓG�*(*ƗT �ҟ]bԊ5
r����?�)����.��o�	�������}�Z��G�/��m����$�T8�`�7�IDr���� ��ï�ُ���H�߾}
|NF���*t+���ِ�"*h���ۻ���kq���7�5Ř��{r;�֜�,>zh�#X7�+�R$K�x�1֟��l�l[� F���j��f`r4��7U��{ܨ]�m�ZL|�$��I���HF�}�?�n��C��e����Ey|z
���Y���4��H���_1�A-;;�sٛ^l�NӁ��������xk*�s`4��"�4���l�E�4�>�g�Ǥ�⪨��` Y��1-�
;���~C����2S����#NU�lid��#�KɄ��́���J����8i`� xƧ�6眄c��2��;�BZYA��yx8���BU�zH��=7�Y�����Fy�}4��T썦�=�F�����g�~n�&�|����@��<�;�O{���I_JYB����EcXKl ���<W��ΪT���8h��RR#��3��ٹ�şk'���l�&c���:��>� f���"�Ӓ&C:��G33�|��C��̦��GGLf��2Y����ٸ�.ԇ��k;;!���k��*H�ȸq����bHMq���N'*��?O�ӔQ�F�:��ϋu%7IHI	�x����H�m�mo+pJk������X�4,���{�B'��w<ݢI|dHEEmv+��+9�Dp&u�Q�8�y�VZ��	ZPJ��Ba?|Ш4P2Gm�
j����c\�l�f3�z�M�����s�ʾ����T��l4����z��N�e�i��5�8�}s�e޾6 �1-��F�
�n�-6��o59��e̋��c`b:��}Ь}AOO���H�%�hl7������'5��R7^�c;;9�d�;AA��yr�����#ůii�%��Rl�CYғ����=�ϲJ�B�vI.�5A�e؈��Y8S�"�HLxbZp����LVI@L}r��y���v�TH����	��X�,>�)Sf�����~�9x��R��;���L�����J�������v�X"�~�hÞ}۷�_[�O��U��m|}}����YP���!��������
x�a^z`����_��h4P�Z��\�-�����L�#		�8g��#Pd�"#���ss��^Ъ+��8����?�=����/�t�X�qqg42$�L�fA�{��t��Ȧ�_�J�缩2Zb�EG��G�{��H.M���7a����B,��Őa|��@(|4.�HO�?�i��m��Rr!��*�ǳ����L����,�>{�_���_XB��#����~//g92ۏ$�y\�A�o�Q�������(��x��3,66ES'99#'e�kR��������g�K��2h�#��ٙ�f�p�A�-6ؒWWU�������%^wAQ��l�6J�"�����K� ����*�}�f��=�Ӗ6�RGl<�ϙ����
r7�؁@����=[��~$9΅�b��r�q����,:N������k��#kv�d��uQ���^�T���bʙ]��������ZZK9_�5��BytkJ�F��o���]E9~�
1%PS��?[k*=��Ȓ�#��A���]��	ʣ�D�R�0	
!��K��5nGZiI開t���a�Z����'+JՒ������PhBB��Aug����q�vsk�H��A/��vo��IV�V����޸�h����IIX�K͘�u�>"�LR�x��&\5�X�6@�ƛ,�,�����.]2����ϑ�ʴfSG�!� �Su��f��K|haY��dnbj
�)��~�I<(�5�f�B:������y�MLf�W������`�k��w�/�­&S̟�V�V7���]���[Հ]���~�[�FRҕ~��+��"ƻ9h���I��������{��bmcs��t�2.# ��t�����)[����zz1�H8��啕���Oo8����}|}��vsX��S3�}�M�����I0����M91c��QNmyIt;��{�����q9OB龲��t[' �����/��j�Y`l�1��R�n�������r��>;�T�D�uF�˚�ʊK�M9_�����#N���š��X�/qe��$�0oYY��cji�j��[{ffT��FGFz@�3ٯ��=C�g�8����i�OSr����xbm������վ���6)''.H���|r���22� I�6��~�SL���v8O:æUg������񵧧'�h /����v�*����D�@II��h*�Sd��XeW�_`�N����+����dZ�ARd08��ui���[�Ϋ������1��d_��l��g��j
���d,@���),���j�~���r��kq���a<LB��4��}��4�{��x�{�nR�AB�éM�o6oS�.̾���� �9+M�����(-9�t3[�;8(QZ�ՠ���-&&��ir�������Z�byy�@�+p6���~��lxı�:Jr��=!(=�W�������۳�I �T):*/������n}wONb76���g�@�~�^�?T?=3u�Vh��焪 ����+*$..Nu��'���y�]].��?�a9[��u��ga'!�jr��ZZ���W���%LKk��?̌����>2��DG���Ì��+��8�[���L$�p;9yX&������������EU}�D��#�P35�޵�w!��anG(/+˃^!��-)z^���%9oO��_�9Yʤef"300��H6|�=���0�C����Lq�����ϼRZ��!� -Ibaa�]-B�[bQ�]M�W1���Uz��ʵ�0БZ.�iNU���	q�������g ��MRR�A� �EjO�.`fv�k�VWITUQH��5�\]���'榧_�E��CW�D��eϟ�sEM�r�.��ͯ�Į�?'L!���q�
��
����S����<6�s��d���)���JP��R��"�F/��_���Lt�TW�`ԣ.{�@M靵��eE�]����IBq�:-�۬v��/�IKK3Y�~�^hC���`�և�����g%���tFFƸ�+P�˓|�m��M�Ύ�n����ga!�=��8h �^�� T�^	���W��2G�!>\5�E�l�[f4'����HKK�J"���' ��d �H�_<����9�bP^�zex�p 
i�� uUe:�U��7�1����"J$���`<�,)2_lX�N��.�8c�ҙ _RQM��Es˫��vϿ��e���G�_v�Py�l���4�)�@����o� �}�g*�<��{e0�K]����x?�j�J��SP��>z��D���!� �o�I�:��-H_���B��d�⹹�9���N,�I#��P�Ԅ	j�ff�`��z�/.��r��KK�����_)��GF"	���L�� 5���� ��d@t����U�������T�ST��{���L��Y��l�_��Yi��}��$�b�,�=�ɉk	�xoO�!] � �.�h"�,��7>�p$��P}Ъ7�����Ri�W�GK_����Si[ί�ˎ�SUQ���Í ����;Չ}S����<<�ٌ��{�ₓ������p�fJ�C��t�Ep��n�,�ʾO��864�H{�o>�� @1L>��$�h~��O��Eb��j ��7�Ǻ��9Ǘ������︃C@@`nwsuen/���:���쎎��X��� "���ED^ �ON�5`�SUU������k��y��k5�������%����"�T��������!��x0K�߅��͛o߿�����G�V8�`��c� @�c�Yr��D�������Vh�D�1����絃�H�΅^���_�n����������������r��h0��#&tyԦ?v/�R<ގ_���4��*�₏.�BerX���cFuoi��Z�%��hã����fJ]�,�>O�|�B��D���2݉�/a�`�~tb��V�@{,���͊
���]�V��G+>g�*J�.���!w�Ġ-��'9t���^���
���1o�K���w��2a�����^���8|waj�a�9?CC�74>%����7�)0W��_���K8�8����!��4��� Xx#@YRO?D'�GFj� �'�/]��Ǜ@}V`�@��L�*���Egz�[�ML��:iz���8��@K���ekԫ��א%՗�'$&B��C�9��0�����Fph(<����0�<*���k�Ц�� 	�t+�g;*F�t[Mjw��	|���#m�*D�"���|�b���Ԕ3j�ha���LCt80��&�!���.��zsB'S�.
{a��ޜ��N��W��u����l^xZ����rS�-W��}�:�.S����sJni�7ox�3s��W��qyd��3�6��ߩ�G��M�n�I�*�_��9��P`%Y�9
E�O�>���ݑ��J�U��~���������y||���g��i�993�y����Mhg����.�T��?�I^{K�,�\�����A�U�@&9�]�~�����Dhq�M�H������o�@/4���<��6+��~	�\QJ'�E`�^\({ 'p;n�"���j�iR.Yr�E����VV����ox�x\Bm����,��
�*5���U����K��pUk�S��L�a�J%%++kA�	������=Y3D�2�~�����F��,�C��]�'�%�����ppw&�i��)�����:=99��*3R֞o1����  LS��[0b�PP��h�q�>�O�m���9FDFBn��`���<r4�������N��2��&�h��j��P��&�N��4�r�����b�Mg��z�o�nZ�Y���\mmm06[^B+ai,�y�#ɧ��A�n!"!a��������B��Pmv������\5���L����zc|���)H���,Q̢�f�N?Y���xz�������wf+�����X��0�KJ'�Z��������D6��l31����,L�z�T:ٖ֙����go;���,2)L{/p�f��w���@#H
�_�խr�z���*" �q��?v������e���)(^@��`������&J�N��VW�$����R(�O�@��I�	\C����J��د�xx��V}o���*X[G@����İ	�*P�7���R,��ǩ�M��EP�Tq�Hu�1DEE_���9D	��1_c\�7�������H{�ITQ6rə/yi�jk�Ȕ.��Ӄc�	�u@��{|d��0n)��a�GK������Y��u��t>��QP�r�3?C@E�Oe��]������j��>E"�� *1o��"������oλr/��{3;Q`P��L>\�;߆֍eF���Zs�.����0���$%�.|��?�6��C�����#(�������Ry�>r��G�<Y�?��ɀN����gR��JRUS� ������;/��+/.Tht�z[su�4��sv~��E�8f��9�G����3[[�1J:xC[�a��Jjj�ƥ���A����}��T� ��7�q�;�]��}��������M"�������Ƿjr�{BE6��0夆�F7sM6K�s�5�����V�$�9�E��R��������f,�����u�v#*���2�r{{�36��B�럩5	�x��v&��o��8�"dP�+�Eq'���*<�p"7��&GFvv�����u�pp@F��|J����d���41##�����ԡ���@")!����v�~��!��^`#�_ ��ӥ�������G�J����B��/6߇��R��$�
��8�� �Ulpa������S�@��I<�nXx,}���}R,Dk��fU�g�_:�F<��|B?���n 3l��,)y`�h ~��Z�cwB>�$##�xB���Y�BBn��!�ue��p�k���
�p�D�###3�ce�����Iȹ����.0�M��:�?{v��nt�zY.nX��VAa��Cgo�l����Ң"8�l�.��ץ.��@��� ��i�����N6�X?mk� )�I陚� `��p�i觥�Elu?��ǜ�ֽ~�62��񂙙٤5v�g�R�k���3`����LM�c��TUg���^�2(|��}F��\YU����V�9���w���o;S��Q҅���O��8�ppX��k�m���r���\P��9�؝�bרc7s��,�(+��i)f�I�1mWYZ�I��^�􎷎�C�E�G|�=-�k"�h��Rmb��Y�*vi6V�Ԕ��r60rNڡt�T���S�g#�-�v��z��ȯ��Kg��F�"����]�+�|�I�:���gY`��*4H�wP��E<o�@���P�y �n�[pk+�X,1
<<<���9��
<H�a�*Ն� �*���<�R��wE�`�}2rrt��?�Y���Gr� bM}��`��c�ڽhڲ�8�f��$7��猆�Ap�n���J�^CQsvI	5��aDs-�H���CZ��(��lu��}\c�Vnꪪ�����qD�Zo���q��AGG�����;g�����N/۝%��YXl.%e+)S���]Ix\�XIYy�=���Sk���F�؜z��-t��`��(US33���| �֏�c���i(Pa��E���V���1�	�c"�oz|A'^"H<��LtZ�Ç����I� $��SG�ƀ�1��T��GXYYada���	��ԗ@�E�R�R���d�ǀ�3���><`Rr��UW�v����W�b���F��[ld�jHjcHKû�:P?9���lrڎ�+�vM�&�R��%&$glx��PK����ef&��2�������5�Fz͟gi��e�n)�_�:�F�h���%��������P�%mR�a�c"��������[��Wt�
Htw*�1��⦦&j��"��o��r�x�� aSY-12�48rb�D��A^�e�����q?���145>�x@e1���� 2�����v8���T��zU/@D���Ĥ�d!
������TT$��'9u,�8��`3þ�+���g�(Rx������La[!�G�d���T�GJkJ�z�����UD^zAQ���(�ۃK)���tMf��䞈�U�o��`u$�����{{�&��'��&ǩ&ME��Ce􊆦�����������mm��]a����4����]��8�'c���C���7T��_�aK�� ���I�������G�a���z U��!��ֳ]%��[�ۭ�)���XW5��2��#�-��;9�.v94��A ���+�[�.���iH	kll�Epגɣ�W<�ܐ5�s�x�RG�Q�rU�Q�S�o�3��^��G�eU1 Suus+e)ۀl���!�춸sK��}�g*+��0,¯ ��W����X�F���X;�WRRs�$�g�Uee�����m�ȧ���ʤ�����Сq��$�v����.`m2y�Q���������{����B�j66l�9����"�!h$1j�ZCL�!�??���|�/?Bo^mC%������������� �[	�1�-111W�IIA������y�e5�ll�>Is=�f�Y!�33d�33r5D�3�m��B����nB��UU}N�5��L��� ׽\�\����PH������g�=��pk\�0a,�<ӄr��|,��8�rS���ÖЕ���6����0����v�!jG��ft��Ly�lR� ��|����yA�f ݒU�UO�eѳyf`c����3�Ʌ	e�h��0P���q�g���� !d444�	%c����JiB��U�qRaI�@/GǏ::=c���3��CLdC�\��D���W�����(���9��J:pgy+�tQ.�EEdn�y�[�$�>�A������˫�j� JI��n~a�m����5-�QAs��4�Z)�R�ZE�Sh�t����z�9߀,�'&j�Z�L}�{��h�$��Ʌ򮰼�,.!�9Rx�*tn14�%�&=
$@u�MQ{{{] �a>�������������11����VV�����Ô��_�|�z �~��	z�"mLJ��Y�[�&(QR�URRZr�d]B��x��0
�83 ,��G��U��G,��SGXɤ�x%$$���9��%&�S�i��|��-5%H$>,�I��*��5	�D	m$��,�-���:�L�M"�R4rKKGVJ��1p#�u����$V]����X� h��`�kl%�HHa�:\��g.,!t����z�����D6�.�tr**8じ>���r�%�S�E���y5����[�#G��B�p���T��FF�;�+ܺ�N/�\�Đҽ��+��aeN��/�4!������I���5��⒦�Y�|�ꊺG�E&���]/��g�f���g_�dXs�G��m0�J�H;L�5c�#��w��jtCy�ht�������VD�h�П?���0887������z*�+-��
��ԆxjIH�<<,%�ŭ�1���2w�*4:ӥ������s���1@��?~�8]{�OAO/��z��U���Rxf&a^M��U�3kBiY���N�@c�C 7�_km���ɛ�:�'�	s����M()�!>:���~ME��*4�w�0o��%4���[=>�M!��y��$����������VNh�%ِ�~jOH��Z��X��V�"spp\-�wa�����Ax���Ǐ=���n���C�H?`�b�88��O`�ƞр.�y���S������������Z��xll�u�	Вp<3V�~ z�����g�>�{�0��f4Ǯ�f%0]#TU����9���ݷz���Z~O[X�^,ļ��l&&ǆ��w���{��9��D�S���@�ftb����\?)� ��g�9�Y�%�+II��333�U�<.���օ67s�������e���?�FFD��W����#��Ņv}��3{a�Dh�,(�H
�����c^Pk�3k�\jJ
���DX�͐r.ڞ��{J��3��hh�-*
955u��a���LBV����������*��o�D@��S@DZ����/H�J)�HK]@���D�[�|����{�T_��=;�3s\A�-�������	Y�2��7����i�u�m&˥S����@p0���i��i��.�b���}|پ�7�S��碀�//g��l�A��t�Uq%qqq-?���_�Ť�I�ʚ���N:��.���,���ꈜy��sZ�p`��(����	��������
%�G# ¬��Z�>}V:FjQ2WTSRz{|+��:�B���.�S���Յ161��B�fC�r�\��3iaeiVZ�`���d5)���]���K����ww�߿��9�\��9M��@�+|O8�U�S�c�D���3P>�3~e�B�h𠀑&މ�ݏ�כ��ԯ��V���¤�8t�w��\�>wY���9��A�$��҉II��+�ӰT�9�F,�5����P{�نP|l��yjƑ<��f�bj%����ϟ���!ԲR����v3Uy���;Y�����ڴ���zi_��p�^s������Ops�|���C������h��uK�n�z�?�x>Q�G���T�N��|��Jk��9'�22� ���Șd�dݣ0��ل�x�W�&�P�\�4N�P���EڔT��~Qņ-ͣ�|�$����lK�4���zT��KN8ͻ(F �,P�ޙ{��lRMO�v�&����������)�_�����5ߢ^�T=A�m�\4��ǃnob4�ay�c�(1ѣ*,s�\L�n�O�۽�΍����U���䊔4�)
-C;�c�P�������9lE��F���QYf��u}�t�N,�?&\�K��^�fG �T�	�[x�Si�������ꦘ�:�B�z���=ŕ��Ieԉ��m�CS��n�°�u�8S�@,]�+<]�$o�=�")"eq__?���P�{���
m�G�{��B���zZ����+kiYU�������}#�RN�0mt��W���%��R�޲nD���) I*���K��״q�[QB����p_�MW�)|3��K
ͫ˓O͒���XK�<�slQ>^^��;y�C���C09��
���Y���/T+Hc&U(_�����*Yz��D�@8���������
e,�Q�]�3Z�/W$�ċ$���dM��j6SA��"[YֻR����sO�莘<��@� �+a��N��5
S��]�&a�궍�dEYVnn��x���	.h�40����W���/��Yi=V��Do�l����ڂ�>�Id��TX��v���
�f�4C�Րݚ����?�����`���V;��7�I�m�y}�=�̱L�����_�����'z?��Sx�3���d���v8C]CA�hK�)�BY�=���7�: n2�^�k+c��B����zaTF��:"���=�Z�A���L�7�߬���[�O��,�f�P&��4��ӕ�M~.ؘ=z3�[�qq��o,O�> ����8�yn��J4]&�'���j������L0�
?���30��E؂�;����A����+���l���v��22h�''%XOʡ�)��&�s����5��*�!"�C��i���'��fo���N@sJ� �ǌv-�f���Lb"(�҉�KR�A����pT꾫%�L�y	��L�ŀ!`PI��y����[D�K��ٹv�]���x.�h��bk�r2�u,U�:2����x���a�L)yy�	XI[�y�=>���m*[.C����\�:����O�>���!�2(���3���s,��vo��а����#K�?��./����g�l̍f�c�{\y0n�ȱ�W��	�<]5��%�8 �5���`."�eE_���N̏_2%!���crL�D YR�99z�m��ʯ{��DB�O:���Z�llү��n���B �f�l4� �9�rs5K%0�y���!�N����
^6�)(M�I.ɽ��-�.?�2{_��X�]3U9ڄ��~ ����|��yҎ)�����G.�����r��|FQѣ����5���h�P5x?^�4�^��S,w�������*�;0�x ���lmRb"l�*��tK/
g�!�+>>Q�2��2<T�����My0���U/Jg�}1��ӓG�/A����,=@@uu���T4+7z]�E��ˋ��.v�Oζ'pH�� �-!L�9�c�	��*��Noΐ�}(����V�֌/O���[2~��#�~C04�ư�.yD�
����Gc��������Jrrr�8��������կ�7���-��Ɍ������D�̪���=y���=N���<aLL^�\�)���� ) 3�/\��U�P��!9��X����������R�(.�,�D�X�P�eOȬ�����,[7����j�@ߛi��〗{�w��n�.��Yw8�j��Lnl���5��瞦��t Mv�e��3owZ�2^�D\��]��9��T����T�N/zBS��Qz,3|���i�J��LPӋ3�?kI!�w��l��̕Nj���2w�@DB?��^붧�`�e�h|��5�Ӓ60A�Y	���$���/���@mK��;S;4�X�is+��'���O�d5����� �h�@��� nj]\]i�jh�^nf3��s���B���[�:����P����������Y�Ε��-��BC����e���D�
'��E�'�E*5�^��#I�O��3��� �dj`n����+�c&Um�����3ZK�P�e����;�����Rbgq�����:�6hK�j�'k�w�{)�������u�A��rQis�x �aY���ɹ0Mp��m�����qo���!���W���3�c���pֶ���Gۊ����9���uk�!�ů0h��2��L�1ڷ������8� ?�&���B�FP4��2t���g�鿅�q̬���������0ٓ���鍻�ل�H�q;ڝX��*qTʎE�|$� a�����QizI��:2F��^M��DOR�9	�O�,^ZT�GU�L�=�g���F�`1��#ps�\��EX�����@���� ��K��,U{˾z���X�b�Y,�;lc�����?�@� �bay���ek2��mll���s��LzciOO��A ��B�����CLR2��ׯ27�24&���[�4P�0T�s�aii	��Q���'����OW����>GA3&������M��<D"(�d������ti�"Z[oF�k�@� 7 �
/T�;��a�ʩ&������R��Ŏ��eD��C#�����!p������-~M�սݝ������7�;�{���3��,āT�VQ�$��o�4��\y���)hi�FFF��x��i>����u.u����T���<�&�2�#��-S��#U
�@��{�A�'���Z�N�6��;f&�󩧿�������R �M ��8K�w���k�°:�b.;;f�����k5�#� W)�� ���.�}�r�sN	Q p"ܱ?�L=KR�w=��,j�r=$C��&� �@�rcQN���w��|5Z�-K�,�c6_aE�����c���ʪU3OИёus{y{���'�movy�{����\���U�~>�U���+B,��$��tA��C$И��ӂ�շuz�N���� A�~w�.,ʲPQ�:����9��dIXoԼ���
..���zz��d�P`����k�QP �_�H�}�ss�jt
�@��8O�N��y?}�1��YW
miNOkutu�G@{�|��Q1ii�U			�-`
��G���N..�[��	ѡ�CCi|��o�x�o���tפ����s�ǀW�Mv��c�z�&бNoS閺�$I������P
=��c �z"B5ŘƲ��23��p4���h�i�`+��m���rl�A08ߑ@��r�aơ�����ˬW�%���n}m�L�K���\���}$ !(6 ��/�y�˂�DIO/����� �mtL�q�f�d��w'..�.P��d�Y��m器���(��RL�k,�+-�W��cAU�)\��;�]Fύ��^:X�\�顺3ҁP��ֽl�p�@W�5I�¶I`�ˎuy��(3mfB[`�JO��r�hE:�Ty<R��6hDs��H5F�V�}i��H�48))��(08:�X]ׄ��Ŧ�S���>	��A���\�$���\�Fv ��5552C�VCa��М��¥S+�7W��3h�(X)
" �m}�����?������H�g�gdi񻉎����Uy|}�q'4Q����t��3oF�dT�����q �1 ��dȑ�{�y���7��HFX.�4���xydJ�CKּ�j+h7���.Glo�*��3J;يtaa���JY�T5�=<~����vr*K����N�=�ij�U���b8ݾZ+=O��p=�1K4�*�n�9P�E�)�����Q�O@@ ���0�Ey�7Q��K-�L�okjj6���^{��������iz�e;�E!�7��`<�����������:BS~��܇6Cy��a������t�)�VQ��\a��k�S'��h��U$�2�db��ޑL�򴎑i�'s"i�'�{y�BC���1�$ʾB���ޜ��h�w�+��������%���B�utl�3 �9���8r�*��
R�=�Y�/ÌB TE���Ⱥ��](�]ڙ۞�7;��S��UJԁX&��p�\�㦷�T�:4���g�T��CW�s����C��;�_��p����kX\��K2��)4��*�P��&&:**R�"pc��w�u����Q�$��pCS�a�V�ommA}�����`�@6^�C�} ��CD����:::��ٙ� 2I<�d��!Ї�?�����}B9<q��"M��k���ԑ!�2�<L��a�_vpAu*9ϭ��{������.���WW�+�o❛�����t�NO"'�V�����~,����?!&�Y�pk{�92_Qc7c�nŘ�Rp8c�a�;]��to�����
	����oT�A���0\��f��3EC��)�x�N�/���2r�̀��f	qX�����d�jL�vޝfϫV���zcr��X�
��q�R���������oX�a�4�m���|��Ó�4O���y��"S������M�$��"jl���ghhdd����|�(��^���U����䊟�����L��E�$� ��ڢ�� x+Zo�tM��Y�Ѻ��effzl��;��@�[�e�KɁݩl%�h�I�����Euw�!���>�	�)hf������öG�l�B�ch�VU6�#���W��z?����w����R�`ڄr/�7Z�.����
�󃥍��Ky�h�6`'�[7���"������F��?��&�Ѯ-6y�����#� ���ʃ��9�VX�Ca ������9��VO/��9�����w�.����-~hhhq}ۢ�9�5��j�ݛ_X8�e���=�r�~|F|���s�
}�TH��sA1�N�'��y����}��T� D�5�f�	1u� �:�F��
@��n(q��?ʌE_wz>�ߛ�q��}޳5�D3}u~�xj0��_�3]�QҖ�i�h�=a�?��Tj(�m��� �Z�2�Ŷ[���j��|�$&��d�WYW��d��6��\RdJf��K�ޜ�������O|cT`g�����7��רE|�Ga{O��i&LM��7��c~���l^i3H�����cά
����ZB�2ct�]�b`1&��JJJX�Ak�I�u1�$�S���h��v9�ަ���,4��v}����~�N&WDJ
� ï���'&������|A8�_��ad5lf.H��L@�>����L��+a����{Dd (�Qwr�Jϟc3!beE���W�<����Y������%����������Z1���#��/@�)�O��f�Ī�!"�����h~~>�V0V.�L�dT��
�8S����=N���m�?�
&0l��4O�A:�Q�Ҫ���g�����qF�g��r�o��9a1�0���(e�#�h��'�ߜw
j&��ރ�H�b��O��A�g�x.?/P��
 q���K5c/HC)Y�l��@���c�� �5b��'��<>;�Jq��7���(삶���7	�;`BB:��:p����w�Fo�M���0E��u0�%�D7	Q�׾jL<!m��n��d��b��pM�+��5A����O��Dށ��|����U������w�AS.�á8O�>���q�������{X��> �h���V��r:K�2PKT[�(�:��ˋB�¯��H�	�l�k����/�P���c��m�y�{�-*�A�����Y]_��8@k}	2s�I"�#"��]�

Uw�--������3��������N���k�S����\�*��R� &Y8P��ll�@?��V1y�ޅ*(Q�2��7�,09d�mi�S��%����>{�p�IZ"�6�ᘄW�񪹢G�'�*��v&`��c��=A8,���Y�4�r$��1�O�HW��:^��wX��~Y����ժ��/7�LÔ3}n�%;�'��R={,{Y����?@�-��Ӿ@�{S"̝�ud�u���ܓ������9y���.h߿i��ե����Z��;�=z��Ԧ;�k����{�=�S1�N�:o���ߨ;�zn��&�"Cu)��Z:t�P�ݰhB�9����4m?��߲�0L0L���p�3�f�����͐���Q�˻�LMª��x��	��!�\mŪ� ��h��� ,Sts�&̜��!�wB*򉊞X:����2Us���3~R�����|4��'���~^�9c'F�M�5)�U͗���McC��4�A߫�w�%�4��HлѲ�ޗޤDG���� �t<�O,>�N�A1݁�u(�|��*,�,�(j�B��[[1��zM��j������;1?���x��^P�&7�6X�n('e���g��vAOo�T���v�B�X�!��G�Ő�\K�
��#;qw6�����`a������0"���YS���w#;]�-�
�bе��=qp-٤��I�y��IG7�߈@9�F��⌰c��g�ZB����xt5=2�����fK l��n>Z��r�͠~]�v�w����E@@G��.W��ݬk�����h�K����׉�(�8x�p���+z ���ޤ�+��I�Y�4,X�E��i��������d�!/��n�`�ㇿ�9r��0��W�E�]�7VX�CCecR5�*���2�hV1K�A�vc�v@Ȏ-7/�ɚ�𑕮 B��Kb����*1��fŲowl��ܛy2�/�9�貇�'�Dxc��$�jf:�������4K��&(w�G��ݻ��.���x�]��n;���֩3�\�>�y���Cb�p����8,�(����6��_��Z��xFGR�F&�9���	A�ܘ�B��S! ZO��hx���� t�������;�ot������:tq{}�؄�� 5�\�X����ץSO�SwFl��7�mYEp��#�����|3��y�܈j���&�Z��4��Nw`m�30g�딈i>���5YU**+KJv�b�`���\��D\��焌�M�`Iվ���8gs����)I,*�C�ٟ�s�r�'��*�����K)q�o.�;�R^������ǅ�1[�ip��g�wZ'+�iە�!|� ���g[�u0E�Z�Ҕ�
�ٷ����2�t'!�utM!]�e2��=>)CC���+��%.�<e����w5n�@7�t�)�����N	T�,(Z�3�~��Cg�ɫ���$0�4����f�o���"�^�ð�X{�C��%Hĸr!"u�9ampJ��;���t/|7��3'�>i����e����jmS�`c�䩳:�jM�ga�#6�t\2pE�����Y�|�Vn��e#�m"E\/���7�d�)�z/�3��o}���f�������E���K����u�H���@���gg��{����!9�4Kos���Z������������N�Y
T.b�?}�2WK�Qm���a�/(s��!%?�U�Y��b�QΜ������@͞)I�;E 2G�v��9�/X����T��,[�*�h�~���mc{.���⢩}'�%��K��\��l� �77W�^��>�������@T���]�����+}��T�R��`�|��C |n�E1VM������)b^�\>�����R�?�ZPF�����U���̀�b���H7�E��U��c�Ht�=8�~qgo���|��4��4}��1�T5&r-]�x��Z��)��YC��b�� �0�)�v3��v��A(`�����i@�O)��o$��S�TW��x�K'�A�H��@�H�JJ�0�Yϗ�4�?�Bϳ�������zM3�J�g*����K��d������&�ߗ���Tv��_EKN~N	�u�	9�T�JJ.�~bߙZ5�~w$���x���D�I	7A�g�ܾ����	q���Q;��a�B�ݕ+�Lx5P
�JX���QdkۖrQd�0}�o���w����R�#u��cq)�#n�t�ze�`( �&�؏�� �U��YJ�7���~o2ߔdY�VS�}��52ب�bp?XI�N���~�O�v��$��0�-;p����%�ܪы_��W	�]8��5T@x��m��{g�m�9.	"|��W��.���˵���Pi=\�@��.i���"d��蓋4��l�|�a0þY�:2�X�Z`��ʢ��l�X������=w������.n\�u�Ȧ;թ��>ܰeh��CYYYM��`��C���iljZ>8`�?ԧ���s�?$��K�1�v���at�	�@��!`��Ѻt�N�K4��&�����-�m���� ��Wԇ�IqW��Kb����\�i`m�KBd59�g�-�)r�犛	k�3ԭ�������]<4�l��z)I�,9��V�וW`�0����2c^?���m�է�|HH� ��m��qV��Q��H[g�C�_������YV���}�ci��@�l���Q@�T��(�h8T�;9='�� Z��p�2�`
�՛�^�$��M���%��x��X)�p��H(�{2��1ni�xM4<���x�T|=���)�Ϲ9��Z�L[񱱱A;�z�R��э�Q�d����8�L���� �FO,\XS~��@�F<�ZDD��_���a�UG�Q+).�<EX��w���2�� %\"�~�?!�zА���ɳ2��rio{F���I��h�pԸ��m�JO���	�M�<����Zh�]�c&3'�z��g������b<_�8$�`1����V�׿�1��2�+��m��\I)(�o�1ҩ�3kW�;�����
�g����r:��3���oͦ���ҙ��33���e���`swR����s��2w�)���ٶ��ҵkk�q�|���
�kb�����4�bK���]�Z~瓯�� O��P]���B�-�B�:,�K��dz��[4�5���)������g������4����������Í!�u�+Uʾ'IFEfa^t�tE���1���;9s:K9U�HF��g
"/�/�a/��=#�o��my��#}���]���pг����K�����+��u�Z����ߜ�aY�m�w��c��=ƑP뺅��~�T��o����T�>����Eg�N��F\~)�5p��*�:(��m+���Ө5�~���#e�i;x�ˮz�Q�?9%D�斌�_j�v��~���J��]
D]�ٙz���ii�$$ϰd�1�yB\�'��ֆ�櫁�����ښ�Y&I��]��@*?'y����b;g���Cd�t���־
7��'xk���3?|�Z�_G+P���Ҕ�wD��ͬ�꺴eX�32�����,��ߊ��7��9��M��5+�i$yՈ���+}	LR����}����$����XY���?��iE��FIL%���%˫�8��(|\����q��6		��m��z���Wn���v�׋�I��`�G�{�G0������]�ϼoB�Js���v�ck����m[{{D5'!��N�'�ú
��U��0� ���W����:��Ņ����(�8���崵�c��V���O��i�dm�k��(�vg���@zu\��.�rY�w�x�4��^�[˛�{�@j�%Ʊ/�����OB#$J�g���Ẹ�вѪ��JM-�U����. ��_�v��!!z�$Onܑ�|d�h���k��K����k��]�?�?`n��=+kF��ZY]�A{
�L�A���6U����ni��t��@�x_/�\mww�˰L�`�|ɘU����3���'�/}e���=�m�/��%���[Ѩ>R]3� ��ή��*������)ѭy	޳��3;��(�}jZZ�Jw�.%�E���`�������R\H��;�$Gߒ	���5O�%� �^q����}�-6�v�t����o�U�3(���"�;����v�D�Tj �W�y��}4^&w�{nM��jv�yZ��1�ۀ���n��Zj}�����e-��f�;�U���\��6�{{�8;}�A�u�;��m������:�or�qKU�5�/�D0�ܽ�(-6�6ʵsUd`k���r{TTT��.���W�����R��A?`��}�-�"ID�� g���L�~�g��ʴ���s��� rB���8�0��.N�!���x�7㱯=��V��	Eš��#ST}���|�������� 9v���j�J>�KN�go�B�mr7�qݿ?2��,���~8��[����53���r1x7	u��R�q�H}��j[��Z���2�?��ہ�n���CY��Վ��V��_�V����%}���VeL��7N�Յ��@�ގ��D݋& ���Lu�����������-�vX��ņ7�?��嘅7ꅙ����P�cb^�~u,�������U�a��Tt�����8T ַ�`n�M������u�����j.:�n�xWP�VC|�mTR���\�����!!�G���Ixa��w�7��p�j���6x3��_J��.�.�VQu��Ì�1�(��<H���������}|�5�R�l9�/fx$ڢ�:�+d^���t�ޒ�������H��}k���O�)6vtڠƳ�Y���rs6���<��R�����k~l�'�����AV�M](��?�Rv%�����r��|,[�6�;ɡRV���؆���1�R����GCC�Z5��ę�Q�ޱ@��ne�$�:Y�(�8���+	�f*�{��Ԣ�"�4@�J�|͒W���)�li��a�d�#��%�+'
�O��A�����0���� W0=ڃ���:����Xg�ݬ"�UਤN��RR(�n{}\��O��l�����\u	X�0����r��������8�̲��5I�v��_f��^�32�ڞ��T�Zh���W}P�|y������M�{�\�9�{-K�h�y��a�SФY�b.�#Ve�����I��4�_����JuJ��:6�����(�m������><v�����˜�������.�����������H"N$�����*���I%������h�v6�ae���d��t�P��>��댨!���������\�e�,��+�`o�bʉn��ԫɟ{[�_�M ���mIj�n�a�;���Q�@�^2��^U�cT��>1EL}c�b3���l�n���ul�����������]ᛂ
 :��'N���ɋw+'/����󇈈5��r����1��)7)�T�����ϻ��0�n..<�{5�_��	�8i�p�>�$�7znt��l߹8ӯ�'����?=/�	m� k�������Ű��h��=]\�s��}g�v:i�y����`g��_����"��*i�-w�qQ�0'?ϔ�)��
{:W�m&�|�Zޗ/��X9�|����HH����Ho|��,��7�%��t����c�+��"�:�������7XM�-�o\M7�7�-C�о���G ��W	�v���d��/� 
�=�w7a�����ڣ��m���93�� sP���W�阘����i�Ƹ�556��]s��m��sV�����N+�����Z�?�b0%��Q�}�h[�ݻ%.. �`�	96s�0�����|X�	He��)�s�D�`����yxx>��h^��Q��5��Y8����k2pe<?_�*����G�6\����x0y���^�2�k����ʞ��Ą�(O��Gzc&���
�ĉ"M���6�׿P��/��3-?���TX~�ݟwQ-��G��G�������Q&6~(e�]I��n9��� ��9"{�:\ޜ M��)e�*.�u�|�\w��gh$%���H���NtYn:�v�]�ڮ�q����O�;�[�_Q�(<��܊oD��(��q<vc'Ӹ���1���w�n��1�l+�Z1��ٍ��(՜ȇ��+�<k����v�gm���֝��'j�u��U�Cg��Y:�`m�l-v��2�nn/���`k4����	~?0`N����+a�Q��
����E��.�����3�cA�W��K���;��}*G�`��5
����<�Ho�O�^�<P���k�Iu�:q�8��{5K�sR��.7�-J:}�(�ⴈ�܅g��,�?FIu_(7Ip��G�������9�m���X�qL�/�v/�P��������'��`��H�x�� )>�bO,�R�T���:J��џ��<߰���Ǘ{�s�7��p�Qq���ڶ}%[��1���$���5Z����.vWk��zEX�r�{���s��^�q�q���ա���yϫX;oF�drE���\��*7]��c5p8x��?~ߢ��y�u�� �����j�� FG^j��0j�1�u{�ww
�ٿq�f;� �^���T�.�(2}{����SN�t�/��bc�&k��z�)��Ŗڮr� �H���;b�o�� u�h#B�(�T��>6�N3a]xa?��#�*�t^� �b��z��nux�]�t�σa�m����҃���Zϊ�{��F}�d����>R���C��Ρ���l�-��:o�{s6e�Hҿk���KI	çddD� <gLL%o��~�ӽ��r��ؤ����55`U�|N��MOk�W�gV���^��Q<*�9��߄��D:�_f**I��|de��5���
��粝�Dũ�֩we���ͨxhG���=G����u _� )~9����Kr6�|���<�+�ZK����En�xN����-a�f˾N�z�������q� Ռj.���}���l�����~�H*�u�=K<��cui�2߾q�dj�����7�P6$U��}�q�UՍ��'�1�/�G""����ī��%��Wg�\7g�\���+3s���	밀i�+>>�U==�Q;ۊ��+�����u9�xa�����n(�q8.m���\�,��,�͊�{�)���8uw/���Z�Z�1��j�������k�ၾi_i戆`X��Ѥ	x�C��=}՛��H��GMCc|����f�{���=�¸������Es���LYڤ����/�����8�ya�D��/�	�$���Y�7󟇦�O�_��Ü{<�߽{_�ki�v�ة��M�o�a�*C�jJ/*��~���W��D����L䵼#y�p��T��<ϻ+L̪�N�[���&�	w��N��_n�+1&�Z� �xi?;N5ŕ/�48T���!�F�k/��Ͳ��f_ 2�zrBq��T|N���,u)�^���2�S5B����v`Li�Imi���1��9S��k�rfx�=�����u��K��(��8��W����ַ�B�i�����窝�Ʌ��m�����;S_y���'Y}�����\�j֍.�������GE�ݬ�.��#��ھ�wXaѹ��Z���]JA�k#�?���ߠ�����H���r{�����/�djq�ǋަ���ٙ*��'��	��ʫV��ey���b3���2��q%/�	OE^G�P��*�qU��LshX��1T�bg^T�FPwf�
Xf�n����s}�=��?�R��iP��=e��Z�t�Ay����r�&��b>Su�Sw�Pܧ��T��V��mA��.�9��TLW�=�9^�z�[1��������!�P�Xb!&j*���F:,���V�H���<.���o���q�~Tjn���w���{�Q>�۴6j~0�{Ӗ�8㩿�����g����{�I���DOg�NQQQ7�p4��&KtW.�V���~�<��n��J�w�n���)�����[�� D��x5��R��>F.;�I�W���޵��]�U\BWO].�/��ffr�v�����whv��\MP������q?�H�,�H�N@�#E�l#�R)2������h-oo����􌛛��ܜ�����r��������Cwww Bpqq� Q��+;:����u&���h��߿�NV�{z��&x��^m7������BC�0��o�B��<o��-k*n��_����WS�-�y_`���;;�i�f��/�]��š�Cs���Lr�p��Y��tF<4��E
����=�͹K��*]'2��ѹ~���Lֵ�/��*����v8\�����/�8,4���Ĳ�S+62��9�z}ɄnNqf+�M�w���?���E��jkW;�F� Ǿ��]i=�E�^,�4�I��r8=�=:�C���N�k�W��?~(e����H�ʊ��Cgÿ���M�*c:h�L�"�����/��^��c��p��P�m__T~�>@����@�"�<��YQ���z{{�?֭���p\$��y��@��o������6���ʹ�D�_�IZ/��5x�;�q7���7[���;��缝Q��[�� ,˹[�)vl�4�T�<-�Ƃ��9D���~�j���m&�#�T���wҘ_>J�,�0� A+�\.�-�E�QdW8���>�6�����S|���w�������a�b��.��oДH昴A��t��JkUJQ00�I�j �S12ʸ��"&.n��#ss�����z�;D#l,_�����V��c�^�I�����B�H��KX���AdVVV�]�MLFF���4D8QOO����M.��+�p,<� ����
Y�j���M��/Φ�]6���fA�g���(3n��H㛢�	�)6��<���# ���I����-H��!�Q���;�J��o�`�Bu�<�o��OK�*�Bh�wc�i�[�^�1�K[���@�?�<�j_0�N�����}�TxoifFAE��s�O��U��*�*��?��,�u{�Fʣ�y˗�!��͚�o�����E�W����_����JT�^���m�Ln[�����vU򄰙rSd�Oi7���z�$�ͩҌM�Z��@o++�<��$����O�99�P�4�$�����H�FI1/m��<&�W�|�|Nu33jZ��@K�k|ttȀP���+x@T^�i9D�P~1"I�\1,X�"�������Y�?�{c�e���u�*��\^ol[�� Qn����
-�P�RC{z�(|��-Ⱦd�aنP�V�
U]KKK�&33Sϔ	a\G];>m@{p����������mkk+���r��P���#1eF�o�A��|��v�1u�u��_��r�I�M�	���s\�m�\�K��d�|�ԵXө��n=�SVQ19�r�%�$�y�(��4�P2tB�Lu���1�ߕ��g�1�;�I���F@�	L����<@:�$�!��a
��%/�=�p��s��'|�D�|����AX���JEY�<P����P_�t�������SN��������xxzj��A۰$FA�-��ON�%��K����Iܿ�9Eх�J� U�5�%p4r���wԊ��}�������!�6�v�x�c��e0k�NV��r2Fu���Gp�@�+f�+(�T�Ԯ���Z~�I�^��KwC��޺�T��`��h8��w��[����Rd��m���ż���7sYX���{�l� ���P�O�$@�r��W<�%) �UT���/ж���~h4�J��>�->|�"E� z&�v
��^�*Y.�����6,��"&43��ݹ��_�ҞA����=`s��%F#��f��E& r��r��X^reZ�F%�.&ov&;�|Qc������}�T��a$�s��Viv�Si����`�niyǱ&���g�{>:
`Z���1.Β e�ht���
|��U�l���D�$���e[�������UK4L���[�����Q�0�оn������\) a��0��4]���K[W���:Rq{2�� �oE���'js�`  c�uDS�:��reۇ��An�Īݚ�O������T�J��0B�	������		utw�+]���9w0S����5gb���A���
y���}�c|dY*�����r�	��4�����OR���~'H]g���&�	��t�/�.kIvN��.��s�U;U���<���~:���&�"����;\��&�44sn�mw��Wn���0v��GIb�����ݝ.� F��l��Q�E���O2E4�R�m������ƌA	'pñ�m��U��OH�X�-LZcY�� c���󤶻��WpBM))		�/���!Y��iiA�FC��)7��2b�!y�
1�@Д�M�D��#�x?b��ܿ��v�о�+}4�j�hl��[�׬�^BO��3�*T C��p�R�d�oOA�
UTT�BDvqK��?���p�T�S���Z؀�5�a��}�"�^�\���<Ȃ�x�o�0��Zo��\$�v�υL����b����B��9AH�l,JSK�J��l�zҨ���MϷ��,QR�R��W��-�x�:Ϊ��O���E/[�9��)�F��;%˺�����P����g����/��f@�g0�7�����F�g�F
ՙ�f*�r�&&T4s4Ԃ�d���� ��BT��C����c�wX�:�<�a���/������!�gtt��^��<
�3)��
>&H��α�3�����#!j�}C����-���/�[A�{|! ֭���Un($o2U�g�m�ͣqK8������Do�>��A ~��E%`�{]�SU[
M����q����@�HW�<C�k����>�@P�V�Nęu�n~!�\)a��wq�m+��Ε�+�I��x?�E��j�ښ�?A�J���gN�ԕ
�G
��x4G�6��[|x8��+����j P�� �iw NB�������YYT��h�!v�PQ<:z`@@@�)��	Xn�A���򭔆>�HUa9�ѹm�A�>�U��7�j�u�W{n����<&))������33D��釧�b@V�T�Y;���&w�Dۭ�g�G��9^��^�D���)Њ���*[�6��!+9?���n����q��~a������n��-�S�hrWb�Hv`ڜ���h�ʰ,��kDA���������iA����n�����o�~���ǁ
�9���k��x��):1!!|Zvuu���	>P�B^�2'sd�����Ex�rs����2�6򞤮�c��7��d�!eg��2�'��b�LҠdz�)�4����1,mz{�↪�T�8Od�{�{}s#���:`maxZuu{��	��E>j���?��"<.g��w�Z$^6�;��&R��G<_��\�2j�<��e4Uz⹴L%����E
������(���E�����x���o
�̂2y1A`�hLJ�,��Ḗ�D�ܚ��ɠ�,�d�ٷAf�@�O�m��u�cz/X::��\��ԋ�ʒ#�����m2|�?G��U�nL�bV������ѡ�m ��\�Z?LW���L}Bn��{ {.+Ȫ2�X]���#��y���Bf��d��(V'��$>��\���VL�z~kk�HL�n�����><����h���.�i��h�`GΒ@��.*k���$��w�IZ^k�-+3l*����s�N����Vv{u�RJ��՟�6���_�m�6��X0Z�O�=*�N��W�~o߼i[\$�c��<yh4&!��˫�e����Y�ԙ����P�9V��wW%:�7Q��2����F�2i��8��d���&��x��P��~Gm�>Y�3�׏�J]�X~w݅p!m�R��'.%b����(<�I��J.�M�U����-7_obɻT�wHG���4��lɰ���F$�9�����۞�U�8iEQ�[��������(�g�����ʬ���v׃�ߐ8�*Ι�F*~��9�}��OD¬���������q����4������H�3����(3���$�э̑��E�sfx��� x�<"K|Pɻ{�9`�����f��AjFF��$A���e��]���������;�wZxNcB��) ��Ջ}=�#��*�����22�]�*�F�ɉ��@@��vgⷉ


`U����qz5`.U�}�@0v���atu��+�3���+`�ZF��u_�N����L�� $HVZ���R�x*����������(�3J�2�~9)ʀ��S��Y�M��� 97b^���?���ט����8f{�۟R�:�����noh�zW�[�]7��ȹO����Z����r_a����Y��]k�H��\�(�T�A˫aυ.��F�hĲ�_��u���>���5*rFM��A(E`{� �y� 6v�����`#�Ĝ�˓�/bj�����D�p��L�
JE��`b�w㷓35���P���O���U
�&��ʸx#�GE��N��֎�N��Cq�����X��k����c�j��[z��)D�_oei�!���uH���¤]��*I�Ж�B^���NNN����D�^/P[:b��]o����2�:������\i�?X?��fA߾}S?�{����Xd9PT�56v��C�O��,�V����H�Utn�����sh ���qs��;��5;����H�?3��w���Qz����<��xY�Di*>��nSA�[
��܊��)-�
�|s½�o��ܸV���ȱBG������C�2��:ܭ��|V=l@�ٴ��H��:L�����*�f+�0T��!�V���	����;�|���ɼ�N..�/_�ק��Z�}�� C�`��߿&�N��*�Oau�xA�ؤ�3��( ��2^�e8�	���ߴ���vQm]]
A�۲W�NwD���| �Y�$���
�3N�?�Z�|�bl�/�A|W�vUU �!�W�)��̮[mݦ��Lv"вN��td|�@��W�gɾ�TX|��2\s�b����3�*7Dyy�}�͵P���*V�S*WU�'��,���jM�t;�ܪ��H����1��V	�_/6�hoo_�a�]�B���[#L��.w,�C^^��n�"�g�-QJJ
l�Y�U6��$��_���P-��kN�hq�:���ǈΠ ����f�	�Dc�p�-k�cR��
#L�/E>�ڗ4�D���$N�� �[��0|W��+/� A��EY]=7��A-����e	�|R�AģPq����د_ �G���������wk��>s��wY:�:8=M��_�0C:*ߩ���n'��n�.7P%;B�Ǡ�H?����H�=����Da�N���(�\#.�QJa������ӳk����:��n6��e���t]ȿt�Z�?�kD��d�XMe�n�N�ldd$�U��@�� �� Ae���X.�su�d�K�q=���Xp��ѽ�.���w���陉�%Z��tF�b�L^߃i꣠����V�jrY:�~e_�pqs�2��ԁ؟[���ZE=8$��v�O���_,wF
z���Mg.#)*��D�w&L!�Y�WCԣ��ѫu	7{wd �~�9�#����*�Kݫ��3� SN$��Z���n��`yi��D�ivoj�g(+ �W��]U��y��Ϗ��,q�U)�>���8�J�t�U~C*o��`c��í⪜o���~
oqq��BH؛H�ft��ͣ>���9�*Ĵ�����e�T7P������_���Ͻ�����U��
������5�?>�(�3o�eT|�Ұ�Q�n�ߔv��W�L�1�K�C(li��|gz�Q&��p˕�ccc�6�8�����1x���^^^p@2v���m��:s��7�����BQٻ��CN�c�:�B~���'�y��"켼=�Ǝ�Pv�^�������>}�葴��8,�-�n��c5T���a����������/��2�ȁ�� �����Ϩ�� �Q=aY2;-�h�+�T���+��o�=Iɠ�p-��M�b�����*��'_�>0�g��5(e�c��ȨX~X�KI����������zץ4
����fy�\��`�����������/��Q-��1©�/�N�˲�ݘ�f��c
v��-������'z��Vf0��ha믋�G�<�x�&G���߅j8��r�E���Ϟ�H��ժt����Xa�6IIɴ��ۛ��[�G�u�zz����G&'o�����@�|��
���oJ��%��f�ss��D�D[tu�����%H�	1vK+�Z��WU�luu��݉�U�����ݝ�?�a��m��t��+�ҍ�|z������#J6�lٚ-�d�̊o�O��,��z�:��	O��e��Y�*yf��'��#{O:\��d�>��1�b�t5*���U�ҟ�����>�Ѱ`OW��'J�C��0���`$t����k�&WE��*��̥`�;*Ku|��PwO�����<��`X����_$�]��9dq�C�Z�������}�Z6t����y?E��-��u�\�nu�ot鳵�;������rdb��}���H�L����0=6��λ3ܒf�hu��6"� �ֻZ�Q����>uT[���ܜ��=R?��NR�
�r��K��:���1����߿Gl��ƛ^e�I���9����lk��u��z�A��+m��z-��ҾA��=�E�6^tu��P��oѩZ���,�v��y���;>���M�>>���I��@[�j��K�NH���$$%e�1o�����U�q��������W��|�*]��ppQ�wjmk^1�{�TU�]��Mɗ_'}�}>B��Q���R�)�	#{������仹��dr!!��Du�ն�H����pxFGFZ� D�K��J�f)}}⠧��%L_���Q�Oq��A������fk�ߔ������w�I�S��j�Yn��"���Ϩ�A����$��h1�� Bi�����>�z6C9�[�CNߔ��D�c,�X^[�8�s �u�@���=����=bUP{���Қ�����/��"��r�3�s�{Z�9:��(�\��sB�I�99햼�I���kx@Z��p�kd����zT�ٓ�/�y ����� ̈KJr�0ܾ��>���˂��?�&�>>vs_�m��IWSN�O���+~�ROʩA�w�{cO�k��|÷�f%�]z�Pb��h_i.
��?�d�m��VMY,,l���Nz/����>�]�:ي�G��[�w��˨�k�DǦU4�/����7�U{<�V��8*]�E�����}f���z�K���A���	����%%� �ŻYtuu��)m'�u��������(9���`7 ͸N73�������\�TS� ����,����������������}p�)55uoo�K��1��&���ȶͣ���H���d�K���8�55�_rrL��g�!��҂�L�(7��P�-��������?�泥�z�,�'X'���-v���/���٭�0{Sj�����{[ӑ�|�	��;�'�w���p6�J�@�*3��_hZ�m��}xzz;-���\E�MF����������i 48ã���*G�kن�뇨��m-�����g���q��gk]I].��6�;D�7�z
�ݕ�](%%�2��Iߴ�D=����6�eN���OG�l�`X����c=Q☯�&7���^�;eVV�I�޺�)������S��vq��Gs��<<��#��VY)i���|����/0��Cѡga�.Q�S����������BEHH;��8�i/k���>}�#oaX,�����(��c b�޾-J[�<��Q��ٻ35b`�MllB�:Sڟ����6(�e�M�@ڀ��$"*�K�@CC�M?��Ҍml.������u,��ddd��J���Fj�`���yph���m�2]g8>+Ƴg���#�5�Q[��Ǒ�XJ*��
�L�)1Ƴ�Pl'wwD�A�_c��fe�����}�b�A2����a�����P�<#=�v���O^%�
�S^*Y���v��B6S�����k{���h˲P�{��Gƫ'G1ǹ�Ƌ
��G*_�d�����\��|�u`@�,`�ZԝYa�u�M�ZZD.��Rֲ�����T��lOt�->��$Ĕ�̭������Ó�2}Ҋ�$�BW��Ɨ�M�nD��U�r3�ka�յ��k� �>3�-f��$�~��މR�0��ֻ,�LD;���u	x�������r7���L�g`(lw~��Ћ�/�� O}��K�l��Ay �䜜G�zuN��Qw�?� ��� ~w���l�G��l,rH������Ύ�2���n� ��t�.B����E�D��tu�z���k��w'dڧ��!��@��_߾����%��Uuu��\7�e�k���,�wG����&�FP����_v�V��x	:���3��V�#b���i��t�`3\����b��;Z=#O=��<���Ѧ7�u����������Ɇ�gv�E����s�2]BH�h�2���Ps~uq����s����?���X�񷝨~H�Zx��@���Y���I���y����L2}}}��qU�%�8�f��sv"{�D2��p����2���_H�Mj�0�Ϻ*
"�	Ϛ)��^���O��^R�~�wp z��E/,<|8��]c;�6X=Jj�vg�l�!hE~:6�A��4����vt�	z"LWZ�@�\��/''')�]蟝M>66F0!�U�/�h��ֻҺ����iyx��+���p{�����ۓ�n��22m �=s��p\l&q���hi�>A�|�{;��5�D��Т�n%�}8
X��K�����<x�Ob�OJ��+))���ՙ� �=N̜���j�l~}5v�:����9���J�80|z�������OT�W!��N�;�[�������a�zsss  ��v=��6��tQ��O��N��Cݓ�Z����k���ǫ��g�el+|A`U]����(TWW�\��ţ�����Kb��7��R��>��O2�}��^>7��z�GECCAAq��Bc�ţ4>g�Q>��h@�\�Q��3c����Ӗ��Naf2��jjjO	���ʤ��龙6DE�%0����b'[Ș _����}��"=�K?q�Hi�```<��F��C�$�ݺ"E��j��4J�������������(h!��4�����\=6��P_�`Ǥ�V��8�4=�y�$����7��S��iC}��Z�$������)8���H w�MILI�8d��"�`�h���]����/&s��Ǖ�<$�z��9N��p0�W����c��͞�Nc���ſ
������*ר�l�W��L��>}�ŕ�J6&���1������Ӕ�����Ο���u�4�4C"#�fj����>q߅�l���3�ب�RA��IP�?����)�^fff�����o_��acg� |l@{�<c	
xA"������p|z��`���]�W*$��\���+�Ya3� �Dvŗ�@+���*���8�� ��1�X3l��:40�����`K���_r�� +9��3 �u.�Ȍ�K �1��?ʹ���$x' f�]�?x�=)GJ�
�ѷ�T �cs%�D�� �LUT*o�q�&����Y�*�@(��G
�\$O#�CP�#X�OF|v?"��*�����y� i! {�K�\��0����Й�(\4[�a����Es磌��W$
��!W8_Qw�\=�|�����0��PTӣY�hggN���L��HE��J�|�
=���I�Q$((���,���D�E��ᧆ�$u?Ƀ@
F��6�ְ���+ / ?���
�8�b �D@\ _�wN�) ��g���`K����gaa�o������:'#���W��}�ޛ��ֿ�<�q��NHH�E 9�F|�ܰU������;�:�Y�"������P5����"&�y���G��Z��	`��0�"؁�D��AQ����R��:�b��@`/�E��#d	�/��f�{E�?Yl��`��<�Yo�]kML�e� �m�2]@Q#�����$]�Ɔ1��)eJ�zπ
ku$T䀟�ك��\�h�Sw!�3��]�j�} ��K�,fik�B���Yb�|,bdr���� �6����0����K���$[u���� ��	$&��9S�ʽ�q8ob66�Ă�"<��byf�H����Pm�65��x��V�_���zaiw��}��^�(�STT�&ow��%��8?Z[[���>c֭~/M��IM^^�i����Ex�&%%�2}���_B�v�V��1���3.ǹ$��IA��:�Ho��<�P��BBĚ��.���**uvwsd��H;�o��Y��*�T��'������o�y|=���aHJI�'��C�~/.^&qN'9�Z�@�"ޞ��5i������pХ:��(����u�6wk^kk��
H8��8aN��l�暞g��S߻w`N�`�_|��Z�݄q�R>>B+���$A��M�܀6��N�g����Uzz�����@�5�ϱ�*�ڽ�=j ,��:�VU�	}�l��X��}��� <���������Le]�G&ff���@$��F�kP}8����\�(�b�P�X�����c��R�=��iF�B +�w1�{s�� �����ǁ|y�����/A�i����/L9����<����������U/���,���i��V�U[�u��NӴ&'�l�<?ۅF~�q*���?�yW1�?SԲ��/j% 0ƨ��O;�T�B5"�;��{���+ׯf)7Kh*���od��^(��k�M���yd��edd��M>ʻ231��\��^�5é�KKK����_d1D	xK�Z�{F����B��[�t\WH��:��{{���CCBK61Qa=���.��,J��8K���t��jdb���/X$�ML~���K��)O�����������{x� �͠�:��S	{01?�z��O� (�������ag��OU���Ĳ���W.�6	���}?��og�x+�����~��0�.�Wes*�Z=O�x��@�������ދ�g#|��o��Ҩ�q	����x����GRY���$/�jk��x��+V; ����I�����V= S��/��G}Ā��Wr���5vS||�,d�)v�#�����8X��t�so�{�ԥ�jbx�����8��� RAZ�e�Ǯ�Z/& ������b����n�w[��|w8�z��g{ۯ*W�,�bZP(�VY����|���������*#c1l|*�vPk������_=�ؙ� �M���K�Y����[hb�Ї�����ְ�,%���''˛��¾��/��T&O^����Ƿ����{����P���
^���Ҳ���n�I2��ƽ˸�; ��Ɔ��Z0� Kiz{������������x[q�k�?|�8���㔊vg�eX#��jȄ�W��a�&�F8�'��]ܶ8v��`���@{@�a�|%���"-80�D`�����%�2�Q�&H_Q�[�~:<��n|sD�wy~H	g�ښ��$M����<̅]�WTT,.�}+RѤ7��y�L�`�a�LAA���і���98��us8�HJ�֖f�1j���|��(����k�+��G�`/�y�������H;�f3�84��^x�#kJ�Pl�B
pעK��=�ޝ�r{ L!dln���$�>�{:���O'3����8}@/�~|��W��ʃ
��m�M����S��]~NIA����'���<����&K�0II��҈"!�D���:ou�/x�S����v����������:~T�|x�޻��D�*,(s�n�"�
sm���m��E\����\���nҨ�9����I����dq�l�몕h�Ru��O�F������v�'s�}No���_e�9���#�˖߅�(��<�о��_�����2w���1HTo�JQ�K�3��1�p�7���~333�nj��Oh������\/c"��*,��)|~ݳj��;]e�nw�հ�׫�?P���  �����������[A �1��.��ݙ�jk������|�]�#}����~K�M�������x�NU����pJ5�\���i݇J@V�9�p�l�D&sZ���f�;C
$D�]bB�)�v�{�Y�t8�p��p�`O����ECCC�y�n!���m%J�[�C�B<�Z嶫��]�	�,�=�GE�>bff�\9<9�:?\�;��W���r�^f
�}T��<X��)bZ=������W�=��ӕ���Fh��L��4��t8����v�$K�gêkj`��QsZM���#�J�/�>�AAW�vy�ɸ㝕��Ѱ�� hHD���1��w7��������=�Q����,�($(���Q,�i��Srq򆹽Ŗ��S��"ے�6�^���W�����4˕������)0���--���e@��d�3��s.�L������1�QI�4��_�r޺&����U]Ĵ������lr^����p�
��6S�ث���E��m7�8��� e���B�77&��T'����;���,r����a����K��狁�C�kV�⇈�m�5I��9��ȁ��Dv`��}�A��m~�~����F�����}5_�m�	�!q�P]�0����@3���II����h�}�,�Eyǋ��D�����k��j���+--�D�������;RdO���')�?ϝ	��?~$�=�d��ZZ(���Y�C'<T��<-%�d�����}��c��
vx7�8�7i���޳����~�P#����`X��AB2��l:9$�6��g�5��b[\7zhz�(n<?�"}K5��.r���W���X`M�����ʊ(k+�׿�'0�2�R�A>��*'W����͎������;�el�X�ۚ`��z�aS�3@D͗\�==Z|�*���!��_m�������R-��~�\	&��L��;�f)�`Lޠ�37=�8��9C%��󣌑;8��s�&�+ه�n�):��q���|���Y�����G�s-b��h�����tz ��������'[�)����+k��t�ÿ47z=)����ٲ�j
�唗�q�O��H�<���
���˰��i�|sN���dC�f��C�hKKYq�6�G�,u� �H�hc?����H��iii)� ���l����+�!�jj����7���o�����(D=z$nn�+jh�	�u� bwVy9ƃGO�ݑ>��p�2�#5�u^�ô���N]}��uH��O�'���Ѥ/�##Q�_ F
�a;:��	3R�;��t�mw��H�NXĳ�� /ه�9��=�w!˳�V�����ǡF4;�;Oc�#��gb�D�%���>FE��������^XV+�F784�ki�8/���X
��t���������x�[B��u�Ȑ��m��������&��I�W���&��}�\��VMŤbmM]�_3�H^��د_��re�%-�}|}�u�Z0D����%��}JME�x����z("D����m���ޮ�&-�M�����Q���<�q�jϗ�>۟aiW�"���=�@	��ɡ����>����|PYU�A4k���S�Q�sL}��~�'ܶo�����k�.���W^k(��{8{"���������5W\7�.����<�)���4�$p#�IT��H���&_}I�#Lx���9������C�O4~"�ɯ;�?a!
z�*��L �������
ӭ����W�E�׵���}��;���*�톘f��ޙ�T��T;�BZ��N����[H�tSޓi���D��Ʉ n+@��Lɹ�����L�G�r[:y}}��_������H��KJ~l�㪷����ȳ�qxYh�����N��74)ED
�mK83�͍&������5Zf$��.�].
��vpz�$N��='�S1��?/.���Mbs8��H.=F�IK���W飛��a6��!�5���U�R���.eV�׉�X��3L��������"""�7@~�	LU�j���&�U�tv�ܵ���h��sA���7���^���;~��Y^[��su�+7�+}w.�'�(����؄
z��K��gwgdc�o6���	C���4i�8\*���}qe\�X�FG?$&��f���t�/w5&���Ƚ ���>�ǃ]��`co�v$2Adp��A=աj�âN�͠����}0�8^��P���%K�"�nu����}���kh���6��_����`E�J�͛�B����Q�f�蹟^�T B8��W�_����0Zz]�ɬ��ƼU򍵭-L�}�����w��:���JD5����\��!�<`�A�dQ B����_ܨ�~U��e�a�},������K\b��������$U�++�0�6���g�R}.�s؞,�� �����_h��r����#�����ˏAl�!�� �[�Hᱥ���ƃ���"222�?#�~f�0벲h�8Ԧ����B���Ɇ%+Ϗ�(aI����iR���7������ag��:i���Mi�ϟ�w`Z����P+�����-B�莎��N[2��yj`:?i*��%ީCJk}��$�J<Z���M|�G.@gz�0NPxxx�P��j�U7?�k2�i|�1!��$u�����ɰ1Icqw�VJ]Λ�FЯ���[ $ⅆ���ӭ�{AAՓ�?Z7��N�׮u$tR'����D8����P�e@	�Pq��rd�ۉ=���:���"v6 �Y�}��A��0���ż�Y�$�P_�+犝��W::���&������'[��)��ʢA������&���9��u�X�� Qx��w�`n�������q���y"�t����/�7�n�`.���n�F�" �3��Sɚ��$��wnV��Z�'A*<�l���D~ �VskG`� �VU��%� &�ʇ����;[v�'��K���f=��q�V�K��4�\Q7|o���S[6��[�'�b�AC�m�@0F��x��A�	,������g+� ����C����w۞T���,���H�E�ݾ�����X��K�����#�*9-�33D���啕�yyԛC
�ϙ�#���P��s�
�ƞ���Ww����juv��+�����
3$��j_�����42��D&���l��yE0�|�vx|;}`	�ǆlg:�ؖ���x\(���c��FJS�x�7�E֑�X�·+��x�ۓ�p�y<#���ߝ��11�i���^]�D�6L��vPI����I��:ޔ�$[07?_�.;Y5s�9''6$���鶛!j�,4��� �e[�T�[�>�����X�����pF��D4�
N�M��mO	#����|�"<�����a��j"ϖ��
�UsdDA���_�B�z r��XCrs��//�HF_z89���*�;�� �_*l-�����41f�g�/�=��[��GU�����=E����3�ħ���m�,5н�������ET������?���?�u,�=Ѐ馀SQJEu��Ů;�Sa�Ïj'�
�<Y^;`�R>�������oO�������M��>~|����_0��Pf�"yw{�>��<�[�>��\0�v���y����.����ON&��Y��~B�J͞dI��/ǁJ"�c��!''GײX%�?Y��uB���ɀ�4�0W
���r�����@ ?zJ�����>�_ F��o����&�rY�of-Oڜ���y�NW(�C%ۏЍ�(� ��!����"	�#��'������H��*��R���(x{��b�}����N����s'\[��}��x@��d_��+;� ��&ڐ�q֏6F�7o$�0���Wc2�I�R��L�R��i빏�ݻ�ЖX�W\̤x�"����xzb7U�6;����2b�_P�cnN߁�{���R�ʑdֵ����n�3X���R�oɃ[����֣ �cbg�F��mSwҒj���������N��,����ף_���! -���Y5.W>�O~ѴuJ���dI%&T�E�z�k��̉���>������-��H�R�}F�KE��R2⥭-X=��|�8�La8�e�l���F
x=|���拯�@�Eҁ���HQ���ܒPa��| �n1���03 ��sW<�0?�u���|r{���6���@0A���%�ӝ>m�����$v3�(��#��>�;}l�g�� 7g��З�a7���r�I�b٦o=<xLMMq�/�.U��R���u��/(Zani���b�v�5&�?�9x�'0ŏ5��:���p�-<[��Xõ��(d0�����_n�[%M�/���6�^�����i}����^���T�[�/s &�� �*kk�����@�\YYu�:��~�Y#��	Z羳{�T}w5���!)Jk!F�^ﹽ���}�u�Cv�և��OH��t(��t�B�οC�n��,f����Ր�45�-Y,�{O�<��p���̵���}Č��$��ű1�����˓m\��o��K燫N�ί�Y��n�'��@����D��>�{�Y�t��2�,,,�}}�樔��g���	x�	��Qn�F�/�C�d<;o0)��.��'�A����4HW6��v��n��JI\Bb��Ã�3�s8$Z�� ��u���l�|� v>���u,O�z<��nzzzic(����&>~O��`�е� ��\�A�]��J��B���_�LB��!GS=����~� RZ��;{{� 4���2#�h�����-<9��OR^���0��ӊ��q¯zE@�^YE� �>�'Z|�)�h�0��=�䥈y�Ã\P�ɉ��:���=l�h��.�P�P�(���a7�*��|zJ�&)���ֽ�Twr�$��ʅ�00����E��}n��j7 ����r�>������>f�y��?��H^�g�p��p������7�o�~���,nK��j 3�aׄ����.���_J�U4H������ք���E�o���P����	Nӆ��w�:0�ϒ��h�0�L���1Z�l`m3J���3U�yȹ��΋J���f;+��xF-xI��|��u�G��GK:�?[[{�xl��?q۶��]�ݕ��,M�Z鍡�G;K�ae�;��� '#���Gw1=�g��V\�@��=�� �mAUww�=26&���|��i0�o��fG++$AAA `�L+ � ?�9L$;�P�Nq�.!!���t+؏��ߜ`Q(���稸�Q
���ཹ
�Q�8����$�	U��g{�����h ��J�4�������G֣�º\EH�4��9%][�[�6� �o�Nr�\��m�zX؏u���/��V�*�9�T�G�������x�c�"���zJ&L��o����Ѿ���]���Bdm�pF#��R��]��w�>��[�0���z?�Z�B�f�}��v�⟖s�M��o��tq���:.6,�vD���7x^Tx� %Ճܣ���i��d�3#"�w��5x�z���*`� ���
p&b�NR �Ϸ��f�ÜJ�����>I�����Yyy�r�,}�]�S
����p1}}bS33�u/V��6�Y~@�A�z���z*"""���8,[s�%��T� �<IK`1�)�\��3��6쭉Rvv�%#J��&�³)���i����)^��n�*�lㄈ��Y:�d݃���(递���v�B#��+��p6����-$�DH�ȯ4�t�	�؄U�E�&��r�p��#�X����D:�91�D�\���+vR�
6�|��j3n���hs�ٓ��Ju�#���O����7�ŇF ��&���$��^��fNeÝ����ň��xw�%�*N����_�d���z�܁��+Dn�cg�qێ��*5 �l��']�AD�k]X0,�^hz�ddd(�
��x�bF=n{�_?&.��:���uʲ"@%"|VCqss*�6t.���%�E�����s�搰�s�
m�P��[ߜ��Pow��m�b�$���Ty�>���E��[������_VT��+-�3E�r$#U����/�tY�?(�|���iok�g����}K��V)ôxI���1�%<`U-|/�~�O�"�|;� wy��9wfy�/)�+���Ҳ}�.�4�E,(����O˨�k_=)�b�x�g�p�0�p��.�;�(�qqqQ�o+���dmk+JeZV�1�ք����5�5>��0����h!�(lU
�u]{�H�e�p����fZ�"����j�Є^� �98��L�onnN�7bǝ��Z[[3���Ӭ��5�B��zpp���]���"<���<3����+�����zc�]r۫3*9F[�II��S�sJ	�t��D�oi'�v*[l�Z�o�_����#�V���F������Cb3nEl<O���nz˻�3S�YC#A�t .��s>>�(�55ܛv{s���a�����՜OF\�Kj�<�y�����x&
m�-Q)��	��1��<b�d(( �(�~%������%'z�Λ������a)�T�r���FG� \��+��rxxH ����s��ȮS�����H�����f�u ��zWVUF2��/����և۬�-������%������N�E�&S��h��H��~D���N�:@#�ł]9�
���YN�n��ͼ3ܚ��nx~��I���߿��`tg�Q�w���� ���5��C�Ǫ�\>�$|�l���w��Q��<iq'UK�m�3S7@�1QW�^YU5h�����`I��r��M����C�6ua�޳�*� �КN�kQ��0(�
��{�J�Õ���{7�1��&@+���
A���{�",|��V�𵫭;��o����9q�*�B2�ФQ�gO5ok��-���M\|�s�P����������D���J�ml'�M�/�����w��u������m#A�Ezc�>��qNNN&���B@@`|{}э��G`�h�
���h*�q�Ӳ(���t��#���,q��#��֐{�<��c~���=%�&�fff&�T�z��hb$��[�[��f�N�L[},L�{�&�54����G`��*|n0�����;�����*��A�2�?��G��]z�my�X��w!��a
�c@�f��Z�����LC(�_�-�31�z�r��6�f��Oh���y����̈́S�%��]�.?U��,�`��*�m�':45���Ą��|ٯ99bA��$�?x*N�r�I��'	O���^F��[ h�*+'G	pJ6�L�;P��=��b�upp0�?���y��eɀB�?!_;X�"M�B[5#�uL[��(�$r{NI�gZ�KMz���cquuM���$�����F��󻊐��b:Υ���j�ٿ�c���{ ��ӏ�:�Ô�?�C<Fդ���y����333��_rrd<v�ޑ�x�x?����B�q�}Um��#i��}��ToOw�w��6���ÑT���^~�G}CC��i��rp0�%��!�v�k�n�0�Ǿ{���/\�d�~ٰ�[���?�l~}�3K�WP��#�LAV����[6��z�yw����@�f	e�nfkG`ߐ5��S`�ti�:$O*#�5Y$DD�I�Ȃg���� x��χ>f�O?'&��!�����M抉�����oMDD�9:�3[mnaA�����D���w̩ɬ�0~k>p`��⍨�,��邞4B�J���l���wS<]AL�����؝Ŗ��o�w9㥩֎���X#+B;��R��p!��Qa��V�q��䔔�_�|A^��}��;w�Ӭ�3�7��=h�����j&�l���߿1@�pii���.�#J
�*e���N�o,1ji����_^=����t�qg�U����o�[�/:���]7�驷/Plll`�\�ԓ�!�w���w������1a5���n��$���Oj���^�2�V����ݎa�������oO)Qbjp��Z�twVJ��x'����8�� ;�ݥ%:UA�'6�R�h���d��b�������`�g�o��������؄�0)%�^l���PJ�jkK��>�JpQS[�5}���-������A����0g<V���M,�A��'��mV�\���lS'�\�Bh(���_�������>��\�4x���RY� ��' �pӨ|�����"�p�0����8�����/W���GҶ�A���<���9Q�����M�Ζ�L-Qɑ�����
��MHH�����_0�pWq�tu5�9�w\h,8N�]ͬ��M���]Ns��y�^>CH����L��EtT�����&y���-���f������{QQQQG ��z�r�л7ӑ���mu����t���	֋��|�:ۿ�;�E��/���	^��d�ʡ�K ��g>/���1B��1�Ks��s����Lݭ��֮u�b�M�Qû(��Ҡ�GUU����ρ,��M��-/�TlА�#�~�	VYs�����ѽ�Q�[���uo�6��4~q&<�[���p�__�IyS-MM)4l��V���Ɠ���C��̉]uu�ع��l#{{�%��߼���[yx�%*]e9d�+��Г4Z
|<!	c"������Z�,,)Fݻnil�r���g~Z6����4r�����G� X�{C�aT�Mj�R�������[�u4��[�{���v�X0���A�4�:}��xC ���ˊ�r�K~�&ff��ۛ�J��^2���jKZ�TEg��7����YS�=����"&D>S�����}��A��C��'�N����@�X�6+�tUW��Ⱥ�^���ރ8�m�ǹ�� �5�o?|����-���z@�#R��e���(�c�D��/0�|�Ԫ����+<2�)�֒CS�����{Ϩ��v]��.���Р�" 9�(�A@��snh�ˀ�&HNJ�HΠ����$g�n���w�{���q��q���gUͷ��<U�s������8Ejck� D~¨.mq�� q�xW\�6����L�`���S�O�K���a �Y���j�L	㠇r!%�w>>��SP�(//�9�$	8}bڕ4��o��h�����~r��ݻw�~�h���'��=<-�f��x����l��p)�o 74��aր��Ҕ���d����*0���c��И��R���n�Ź�\��Щ%(����xʂ��̣DԤ`pn+��#ww�z��C!���k�o,�|}����dGY1��M�SС�[��� L�ruk��UAS%��˗7X�M���"$ۇ�*e��9�⬎kz�SS��{')&�1W�͇O"�l�Xt��7l%�@�G/0����T�h�Cb����"�m��v��
�=�,M>�*W���q ��tr�Bu f�j�L��Z����ʊ,j1/o�`��	b �s��3P�LWL�{�̸���T;Ϝ��U�|QS-�Nf���0���p&!)���ϸL $@�j�7n�x���R_�����?7J�Sœ8 .i4����(�X3�ì�z���ă��ZN�I�Z���7�$�ZFUSﭮ� j��u|Җ߯TSW@,]4pʍ���6F����PD��X���0��*Wh�1�ɻ�߿��'dg���f����m-I��)�!�����b��	���Y�7juXxP[f���>�GGO�u#8L�#�H�[l灓4^�P�. <�30�:�t�o߮����`_�vz�A��lcs��������RRR�9��o�܅��
����Fz�U���3������3���В�L��Լ��A�5ee|��i�����\q㺧H�S8��m�� Z�dnr��tv����op0^%[+E�(�Y$��dY��?撥� �Nz��9���|	tX�=Jt�z�+~ ��߿�gW>D��pQFF����˸�,�V�kv�΃�(��
���@�5��@?�*V��YZ7ˡ-=��G�7n���`�x�ͷ��}}�}}}�oWnuF'Gu�������w���s��e��ͦ�t�ϕ��<��{x	���fkk��O��>/��gn�7.�m�� ����c��9����B�w����U��A�C���56h 0�Ct:0=k��(u�o?F��D��u5�k�S�s��}�Rؚٸǭ^��cW�'xl��ډ����]Աb�k}G~��w�Z�o4�ih��F�F�ݚi�.�6,�vg���{��9�*�?�(��DP(��f�lU�G�z�t��aN���z�|�]W���u["8VG9c�=U���zz��r�߿o�H�\"c��p�y\`��ƅ�B��=�æ��A�P�`5nw&-�ڢXuzbq������e=Q�4>!a���row7	���{�Mou��*B����=V�{: c��zGX��P�AU;FEI��ot��x�ta<-=�w���~?�^9�PE[�y�XO�n�W��4���5J	o��Ni�?<\9�C�jM�L-^�ܿ�k]��X\�9���&����TE��x��DP쁞�H����^F�&����m�y*�V�����|�ʘǨ�>����
����v%)r�������1A� @V�ri�\R���Y/,p�q���G�������� ��bݭ���i�/=9L��UV
�RW�/,��n�w���Qҋ�� �x��BϷ�3��66��F��*���mmm���
	��d���b��f�����;�ݓ����Y�jν��D�|��i��/�e�	:U1�>C-o|���a��d<�ƣ:fW���B�""륂^J�
@���&�ũ&+@	&��z�l+5�+����;�
��x*D}�T{�U��(�+HGٮ߱S6�~�r�ʃ)fL��fuc*�/pp�W��ϊ2�Wōj>^Y��t�^�::427o��rg}}@�%����V>����)���y�����B��6�u�ɮ�M�O�sss�~�}N�-�24��&�����*=Y}��� <U:��|o��nm�yM�hC6�p�!���#�r�[�Xb;� �&�J�c�J���z�3�/q	yyy*y�����������*����#�h�����Ǎv� u�
��q/���*�RC�aLx���nCA�V��Lt�!���TKG���GM�k����.Ȏ�.����z���l/�Oe�� ��> �.���di;�`��P�Y�,z ���@@W-$x�!=��r��r���$�
6�C_]~_���9���M���t��!��#	�Ċ
���S�+��Cԥ��A:�IQ���`�-�*]����$IGv��1V�lk��F`T�q��^jZ�sJם��%?%��m�EI+�p��!�js��O=��_[����SS  �d���t=�*vU�����]��pw�v{����γR����!D�f��at�.�&�Qzv/G�FPWo�!�}?�'K32�uo�e���LuEI	$�su���6C�\ 2�F �X-G�QW,J�B2bu�ڞ��O�޽�6��t�jP�XS�e� %Z��V_@e�G�ׯc�V-E�,�B���d*ףWh �b�N+d�2k�]Ps�������0������V����2����p_h�a CV�=zff�A�k�� �ꭎש�Su!����~��u�:���h`�P��'�� I�0�r7K�=��f���)�v�r� [�baa!H�m���' T�Z[���3j�P"4$$$E����.ƨ��Lƒ�8��Or��!�$?F7��1���h�K��N�www�g�>|��Ƭ��|FU��C���#\���.}^q�ਡb{$R�i.�}S�y\�M���o��W��@����S�)d2]gª���y���Ζ�K���r�(�,ι�T�1á����хs��B�9�Rn�S:N����mg�]7�%�={v���_��B-�\�R�Ϣ�!3�,S���$����AC7��g��5��H\/u9� g�K��g�Yof�v�bh�"at�ݜQ�����g�R�`�7s�jd�(��*�����\���:&]VP�?bl���::.��Z�1��6�R� �1��b�F.�$�M5(�h�ǎ�#ՀHk�l�D��w�m+ό���f��Rw�3%�� �x�S��i7��B�7ߕj�'9�r��[�-��I������L{2x�6��yBS�\H��{J��}���@���q%/�
�C~{�<\E��}�W빛����Mv�K�[�t�a�h4&ʦ���[L��&.���'is�ۦ�ީ&�4�}��Diz���������[ ֹ�qa���í����L]i))YU�{�S��2K<���4�G��A �d�����
n�t�w�L�(�6�`;��{zz��lU+�kh�� >������E *�� 9��-���b����YR�D�����e/8���ܲq�����:h�Vnj��{rXs�;�T��i�s�<R��VO�D�_W����H�#���C��o�|p�r�z����8�՝	4&M9�u�\p!#Og�g���<`PUOL�������,��v� ��7����M�ʻ��a�҇�e�����u������������<�MS6�� O@���D����)���̕;:��ri �p �'>3s�+��R�2�wCz� 0Y�U�l���X��* }�hy/�%c�{Vs�.� �ٮ�7����ڄ� �+�ƺ��&r0�|�33 ��,�X�.�hyFDD�4^�ٛ��=<�ū�`w}b�S�?CW�ioM�B�m-H�T31(�`c�y�X?��TSg��o�����NW��M5A��WW�D��?�/-����{�Owb6�w��G�] : ��kiQ��wt\��}h���� T-`��Z�i�֪y�4聴�w�.ԗ�<Fff> Z�dg�!{�fW܄^	�o�FMY�$9���E7��N�@utt���qqq��cbb2i"$$$��ШD�I���{w2H���02�#��jjj��*yv�I��)�o,���_ ȓy+�"�
�������}�`S@M<>V���V̏��W�!fpd��{.!Hgoc��S-����$� e��ꪕb� �������и�T��	'�4Sm��`�n�@Q��~�l,�b��/�OpP�T̆K9���� �Z�рu��>?~̘`��ѧ�����"��RogC`����U�����Q\����e�`
\�+��pZ�8�r+�~����
�FΧ��:2k9��p���_uu[��2)'����
�mB�{Zj�'�z�����<����sP�X �&�7BS��Q��)))�0�z;�������E��pom�7��z0��565A/����de	Zi����C��CM�(� h#KK!��0i.;8������ːa��p,y��S"���C�1ݥm/�ܟS6j�'�a�M���)t�	
�ho�bu	���W��}?neq�k�/����7�l^g&k�/'�I+���Ͼ�`�?ج��fQEZi
�-�����/�t>�P���߼Ғ�<Řc�2�������O�Lur��M�<Ų��32\��ƾYlO���nu���C~�RH��N���P�C�CZ�>i�-j����#�\�hR�t���J|K�"W���ϟk?�6{20E��n�Vem�_����RW;�ߐ�*.�*�����]ɖD��rf"�6�-x�"ig ���2��XL���M�-�)Ԍ��$���@N:g�>�C���BM�����f1����p>h�3H&,񹨫����p#U5w11#��Lo��0h8��[;�Aq��8Zh���Ό7��ך�9��4���ks�_��D5*��o�P.CG����X^�p�ni7��.��O��*�m_���f,k�l��O�@�{/������ὴ���~6�����⽚����OZ��Ri���&.�l��Q�l��| ��D��,��m��qW�6�%�.�qً��+ �PXOE���e|�=Uy��Њ�f��c5����qH�O�gy~��&�T��VB�F�m��ړ�.S]�u��<��/����glJ����|�u$ȵߥ;��Ö�w�x���9Ẃ.�SM�.���Gؓ���ɫ����q��W3��d��XW��ϸ@v<������X�g/�\�\1�qi��N.'<
���Ȱk���3R�r[N=��~8�a����mv�L�j�g�I���c;ǽ �v4��\W(�ۜ��z|5(�Db/�b4�%�-���:(�̋����Øk�-ZI���(�f:Ɩň�cA2~��4о��M�%Q����1�����$�z�S�.�����9#��Ҷn����F/�;&ޭO���?_Ӧ,�k�(��߅�۪]:j�?e�^�z	桤?��@L�o����n������w���@m2�S�4_m�3l~t	M��=���#�q�E/���u|���t�D�$�B�sR���
&����nR��?z��B=�z�S��c��t^h������s�C䑯.�hV����"#k$(�oFXW[]*�o,I�\ ��O����px Q���^�����>?55ł��cfF�8>�4��G�x)!�|%�� 1�HCN��"�~��@O�buh�>H_z�����m��dS���Y�<ݙʧ*��i�4�x�=�\o���a�m�����p2 2tk�� ���Oɘ�!xU\��G��xn��&�[��0�[9Ÿ�A�%�p� �L�!r�8��ˌ�K9��1��{*��C󖓃VѰ�z��w8 I�]\A�E�� =�l�i�XO�4D#Y~�E=�v��a���D����A������XG��y��ՋV|�#�	���88(���6�Wǥ�^ �|)9D;�Hc����mU��uR&�IDέ�\&�캎�y��C���nwd\N*Gwx6r/���"���r�v���0�M����2.Vp�|������֓����;j=�9 .�Pf��":��Ãy�՘K����3S*�����=,�{��;�[?M$�ZK�]���vQ��s\��DLO�f�wV�>%�{d�3w���V�$C�����R2����64SU����h���LDV���FL������V�&�ީ�&�F�]��,1��o��B�s�(x0Fh��"88ZF�of��{Zr����J*z��J�k��=D %��ܛ}7������6�� �)������@��V�6�da�Kj��B\{?[��9�;�K�3nA��[ ����f�z��d�G�D���Ϩ�S4#�h������ >o��mk�G���� z2��β�mws�璼�-2���Y���w��
M�H��:�C ����Ȩ&�增B����^ I ���p���貽姯�s6GDF��A�A^��v̞���@F!*<kEX��T$�6FI���"�h�BD0ߎ�E��L��W�� 9XXxm�4���=�7!��Eg�)p.4����SMu��zsA�	��ܧ� ^�G��/h=-������%��	��iq@���Т����h��=����sfT�ap�6[���޾3x����>2Z��-@�F+�-��/�Q�����O����O�=�ۮ]���z/1�u��}�#�GL0�/�`n�c��b����sC�����#G]鶺9��~�Sp,m�1g�� �	�,��A2>w�a(V�B�]�r��٬�ɢ�;9K/Ο�_𚔒��L�'���a�|�ˣ`��8����j��.������wݚI`5Ŷ�*�w��K�166��d\��ȉ���w����+i���o�j��5P��=��\�1ET^�I Q��L��v������x1r�e~��c+�:F�hM�0���S,IK�UسGܱ!����wH��~��1]���t@izC�U8�2�5���'�(����A�P�������n�> ��h��k����Ԏw���]�u9�KI.!����mr�q����:�hr�EՁ���W3� �G�K�t�'��0<)΂��k/���ݒPq9k�^�q��%�L�EV�n0�j;�oe#V7ݎƹ����c�S����64DL�T��z�1B~a �fP�����;�����FP����0l�
͆o���֩RP�V�,Yo$��öu�e��I�\���{�~��.L'�K�B��	�v�T'ʩ|_3�<'.��[�_�����fx�S�1�,D�ٳ��hW��PI�"E�ׇ����g�6U��uuJ��,(�Z�����)��J��1(j�sU/�Y�\�}��>0p����H����(���a�}a�o��^~�6i�,M�+����1Co��'��}^<�Fw�!mKmME�
gM�;�֍�`�7�����q}Q��p�[����#�2���}]�ː��(qÏ���b�k�����d�J�_�W�#@B�Ǯc.�b|D��Q�?�ê�u��s3��W��p����d��+C���b�y3o��u�Yr�&�a�~ȓ�h<*����Qe˻�U�T��WxX�㶟,�����N�$^��n|�T��kB~>;T �����=�YM]D�����xFZV�@�F�����������rD�~S~�h}���C��NH:tJs�AoU��D�b� #��m��$�栭8����, ��t�!����@zϜ�d̬�b|���ȤB��P�5���ü-�(�WS�o&0������\�壢A'\1�m�zaY�Ȉ�꾘�g���R��7���z�
�hk'���2���7��#9,��"/A7>&S�b0��m�%*/��7���������,��ƶ��2	].�[#�y�'�4�@�9��_Zm,��"�����+6�1����08���`���8�\g~�s��6�K��
5�MN���r��W�uu/Tjf���x����бs}�Jޑ��cDlQ_�hd��n�;�
�����K5���E�����:յ���j�G�����6��p�<"�lC��z���C4K[�}�3���buLQ�醎�9$�������>� �%��c]1Z�H�zh;Z_`���p���i�� ��B�j������Z�8n����bMR�bo\ �%�1����M��������+E�3�b�KIa��|�q�����&��r��#��4j�~���;���Mj�PL�;z�E����B�}���Ts��ه�Z���/����]�ۚb\�UM��R����u�W����]��%�=����um�职v���w�b} N�,�r�	�]�n�%�z��<..���Q*���ő��M[�h�bdf"�?2�)�2���v�M���ə��b0��\�h�oF���M�,���Y�����"xv��s�1�J��=_u]\}���v�"�r��5��e�{~����B� ��G(����uP�ʁz��y2V�X�k���Kp��Y�5̑LBp��l=�e�AQ�W����d]���+v�$��T͍3\b"�3���}$|��I��{���ߑ�v�|��>+��#��?������5���xqqIO��{�Kyy"h�s~~_��% N�} rr�ZZ�}���A���	6�4�>�aΐ�=���P��S��mtBK��[K�����u�=��9z8�ҳ�H�S��^g�1Y���s�����{�{��S�R�kiży��z���d�l}���L�-��kQh�OQV�ڤV-0Qn���H �~���͡VP��B�������� ��wBT�v*T��h���fѐ���HWw���r7��h{{@cԈ���H�I��r�|��
���ߚw�����5'&&��3100H,���J*|�-���x��M��ބ������-��ο��6;A����}�
�M-��\�b�F�}��PP>?K��v&��k�=ۿ����@�,�C�{���5l{Lp�p{+s5��H6v��.4�Q��ۻ�+X�4��fp�٧�e�_��d�6��H��Z��x-��ѯBd���M��RL��.sR#[?�ѵ�C5~�x����7~�m����tq��4��fB��l��c�%o���e�H�[��c���
;��ѫaۖ�vS�g� ���d�:�F�c��\
����w�m�~h���$��h}a���6.�s.J�����f;J��@�ڠ5j7d�����u��_�~Ř�� �|\��MQSC9j����lmm�+�pN�jW �>��Q~6�����w����D�***�ؗ�(M��x�t���ϼ�����g�@Ob���O\\�(��8��'đH$`v{��8k���?t�:�;��N*���j��6۷B�� w�5zv�tW-讅��3_Fmr�@E���|��SVSw727G�*�״�P��<^��Q��[+��1j1����U�m�!� ��9d���v���_7���g�ZR����Wo�y�'� \u&��}$��g��
h�ν{���uw~�4M���nc���>�ò�5���ђڪQ�����2��j!mh�͜�:��30�NGRW����	�ѝ*Һ	���/b��ϧ���ee��V����3��,Ay���9��m\���O z�~/�PX�I*{n�� �Nq�G4���2�hvV�F)��}����U����||.<��}'�B\]Zn�zinn�w�{�꿰�67�JrG�g%���S�t���_rr�g�O>u�������~��2?P��n_R��a"��3m������)�ۭ ����S��F|2�g@�'���@$VPA~�]�BRT�{��)���<�O�;����B��� mI#�H��'-��[���xo{;�d `ƿ��^[�3� �b[�88RE v��߆ )�;�5�zg�E�3��=T@\��T�p���2��y��~�����WM�K������e�wQ��q=�#ץ����=�+�)�O�܆�Y.���/S��I��_�9؃Y���>�Hd� )�'�Р��$[%�ޗ��,p4�W��G��5��z�˷t\�+ �m���ѫ�yU^�7k?��z��&�0����H+H�ko�N�ݝ���W�1����М���1���K#���!->�=��*��e�oE���Q���oƃo�\���W��dh�Tk��������[�HٽX,�Ve��d�.���!e��[Rn۸�iD>�xeC�#^�7?��'��+�Y�4me�궀�q��9����y�8�!�	_�f̆CUVV�N?���6n^�r�_�m��Zz9W|�YŊ��a �Iv�xY�x�t��y=rԧSVH��g&*�U���M����W����v٨(�P��m��τ��3З�rl�OH�������-4؃�*�9y�� ��o��f6���[VN��30���T�UG�lm�F#�z�D.㤡X�N�����f�/��	�퀿�C��r��pi�J]�[e<f��`5�Ewк^�6wN���X�j�YuI]
��Z�WI�S~�
�������{�65�u�,�73�{�A���Y�,�|Ư%��w�a0����o@I�<:
�����^���D��.��oÝ�yݟ��g}��$�������g���0��:gb=d�������y����n���ģo��T�HC�_P�1�$� D��j:��K@_�;��r�:O��8ﮝx�����<��A�1�rЖpr��C����c[
?�j���?�H�]���?*��݂����e7w�d+��QPxr���:w"j���ʍ��M�X�� ���J^�m�B{�t��-��z��΅6M������=��f�'�r���.�`�?��� )����j<���>WG�mji��Е{�g�x�H�!�wp+n���)II
�����f	����+δ@!K���@�[,]omj#.�ޜ����'��{ 15k��
r��� �� �4T��1���~�&�\\���C�pq��m�;!��*�V2˶��t�?2A�<���pU�p�/�M�ސ�Y[D�:lm��{�H��/(�X��� ��S i���0iF�1�׌f���;���=6�EW��eE�f5;;{�Ī�tL����squE�C�U)���e��9��g�@{�4�ы�7���ܵx��ޭwI�0�\|q%%�.��ܰ�p{�H�|3�Ut����3�`u������eA�q@��΁���F0�3�;�Z��bU6�8�x�X,�y���#,	�}s[��y���4��ت&���@�_�#�?\"����Ji��nk
��m�>�9�R�cC�i'��3qNF$���_��AN�J�>���%G�ނ;ϖ>�j�r��=bM���@���E���� N���	J4$?����ߝJ�Ȉ�U�?QM��տ��/ky�O���������9H����ҩO^Nl?I�y�|����k���=�1�;u�6�8�����_�0�
�[����k$`��f��Z�y�_���ZcE��Q ���f���{PT��~�2���=�2E3��ؿ��4�v����Zn��f%�Bήڵ����,Gg'��nz��(�������1���bi�U\��(Z�;��l
��=&��rg����C�`0c�"�%�T̠���s���N��s�e\��(c�\�=��C�X_��HJ�?Wp�;/3T�P�Y�|�ፍ��V��Gr�O��GG� �F#^��4�?c]s�K0�����e��}�9$�:'�Ő�=�bS��a��a������+@ �^��Q�Z�uJ[�*�9G�qM{�Qe��( Y��z��'���%��0r�r�z_�^qO��/ *����-!���	$` �� Z?�/Gr��|B����+	, ���,�-!
P:��]�� ���n� ?�C.K��j�#|\���CŐ��Ǿ���_I���ۼ�fQ,+5 k�#�To�ť�/
�[Q%<��/��|2�z}���x�w�ȅ ���p��L5�v��(F��X�~ "�>�cn��?ɛi�.ʹCR`d+����PB�J� �$�����L�^�h5���q����5��c��)`Bg�/ީ<�2G�p�O�k�M 7 �7���Q�s���;�C��1��)AW�ߵ�/i���e�]g��#�W��{q		46%Co!��� �����[���z����=���� ������w��s�C�<�z���<�;A�剸�(qq�l�-����;�"|ډ=]w���)>��V/�Ò�Vt5Am�F̊^�	H�����UTྦྷ�t ����U֌�Giii���Q\��C�P�(���R�qC���XCӫ T��, ��RRMo���|nhhQmee �� 4���X�.�~���X��P��'tZ��aL�Y��GO�8ΞSӗ���*���d�I�Ę�M;p3Ԧ �ia�>R�3ғȤl���tȿ�Q�_oh��Z�ŌRU8���|`8���(@�^�c[�E!�F�G�Tbru��2\��cc�8�v��Y\�!7ò�_����rcV��U��ix;�����Tpqq�����-���)���yOPH�hjF?��?G�������]9��H��	
�ڱ����������z�*�T���pp����|<E��Ԩ�����:RN�'��b�&FF����cVKl�g��A-�Z�:�|�������$�K7}R�G�X��н�'9��ݿv����<����
�j�*�rYW*�����$�"/0�<���������4b�q:ܝ��r\���A-{����AG��M�y":������r�U�ʖy�)��j�vj���>�>$&��}��}��I�/Y=t����+&<n͎�2�mt��{1�uHҦJ�2�Z�ra�Κ�uӊ��߰�S{9@����u�V�1I�=F%+��\m	g��]&�vգs|~+�ܻ'���v���-�;����9�x�	3'�	ޱ,�/_��N�G�0��\�i�D��:�^_��~�cL*9r�B��`�EJo.��gZ����"�>�z~<Ѷ-�u���f�WD�����(�:���ʐ���>I"���-0<*t<w�l���3=*�E'��W��S:݂��c�;���ה���͑�qw�mع�	O�M,ֶ�ٜhH�P��Y�x};�~���G,��S�;�^UqZN���K���Ow��p�i�29�9�X*Q��%�=j�&w�Er^���n0ʢR�d_�0�V�$)d��3���0(���1=W�j�:b!0���>$kSG�B� �_O�h��Eg�$�f��+e�ڱS7�	����ñ��i.@
T6��۫����FNg�V��.j���)0i�`���N@>?�|��%c�����)n���,��z�������j2%�qޘ[~o������Ka�9p�U1G���iJ�1;��~n�ݱ���	�9Ǭ����޲��4b.���EEE�{E��&��,ٗI���Ƕ�����,G+of���i�o��J)����G��>���&ȹ���6S�7n/�Q����c��t.]�C$�}�S�D)�耀���!���r�칋����Y���f�x6x�2++�$s"޿ם*!eQ���'�/̝ �N����o���< O%�`Ri^BV���Mk6'V����$+����pS�D�;d[��`x �����<�+�f� F�Wy]�����ɝ�U���ɾ��2#�8�+�MK��~�p�Х!���GH������M� ����M���fY'Ê���&�}?��6-;[�����.��PR��e5�ع����̹� �)={��)va}���q�`�_���X2����5��d>�%L�`����cQhh#��[�F767��(�������Q4Ȉ�Ԑ�9�� ���K�����~s�?JW[��I�`��:]ش�	ȥ%&V��z^�H��H��h#rmx��y]�(�Ә��VB0�*�ر���6��N~��:A�����@6;�k ��G&ʷK�"
��tﴰw�ܟ�Q��`?^���E���"�4��*^n�|'ѵx�t���L�N�������������gN`�1��k�W\)66������*�r��/k�it���H����=5�_�ߟ1�1j4וi����H|������'��ƙsrd�7Q�Z���&-%�1(YW'�8]q�4�^#�)@l6C���T�!#c���6���#���N3�mII�E����R��c5�39���m:����y��H�7@Z�@� �Л]���?���20¯hIc�T�1(� >��#���{Gm�Gv�x�v�}{�p'�b�J��'�n�d�JB��C�Hp��X^���LMKc���}$�����_��8�5����?���+Wrw����ҐR(�T��|�RI������hx�y����� ���R"�[C������r���[Ԁ<����TI�t�	(�@s|���=Dqv�����ǉ�?A#��(ݿf��X|���!�� I�]�I�SXs�?��S�e	��"K.�)�N �v���Q��FHS]QԨқЛ��K 'o�@�n#��ebjJr�C��ų����Yu4�Xm
�UJ ��&R'��nkg�� B��
,![��wf����e�b�z�|�|}5<��
_��+pt���a����%���������u�rE.\�xOnyU`,�G�����E�N[[ۗ��<W;��68E�$�Zߵ��F����jlm�_���i�d�nм(5?��.�s��0�{c�S=�c��;� 1 o����%��_��Ҋ��u�%��;W��x�B�e�{o�S���wX��@T�T���PI��+7�KMMM����&��\�@8j��ZΫ���vĵ���C�]�k��@�iV�X�˖Z^�������񨋰���w��Q�+���j�������E�Ͱ�ߒ���e����r������ƣg�׬0	Y�)�P���]�{���§5QKI�����{�Unn�v��N�⛓A�����YY����oO�\�Y���b'�r^kH����ic��H�tk))>_��~���P���4�L�?�CHf��6e��~���P��`�lII	HJ?��ץſ߅��T��D��G�J _��A�-���'������r8H^��%���Ḙ���0��_f���=}}�׏w�Wh�gFTT0Z5�k�-N#�R��������ư�O��1d�������rL�S,�l�#Ժ�Y����~r�����V�ٰF���@�SW)����N�b�ן� < YNZZ:��iQ*����x�����ίr��W���*����q�����]7��CB"�����^��x%�w�|��~e$s�Y�$c{�����ͨ�5����"�������y0�Wy�W<#zRi7z�!j*Y��2��U�	)͚2��X�nSYsS�p�g�+�N{w�p�5�>ug@^U5����%����3�Q�sll6���@`���Au�
eۙV�MGH'4�@'����h����1�< j�n\��x ��U�k��7��.rZ�\���ߝrZk�UH�I��Lbk��y��nQR��wt��h���w����a*��G~�ü9��t!��,�ä�N}�=�K�k��9���[B��'�x͛�M{1j����I�nf�e��
�d�i�A*�~�83f}k�r���B��-##����`Ձ*]W��g��F-6y�SeS-p;r�g������������7��,�@3u�֧`歡ڮ�lX~E��fg��DW�:Wpp�qw��Y"�R�@*&��4�Xq���׋W�)) ������:��F��h��@��ş&�Jۭ|+�������W���^Ul��^U:�ܾ}����V`paJ��`��U��G&��������Z��Y�uK�D�Va3�u��*�A%@gh�J!>$/|m�ߦl�ݻPh�R��j���ω����G���₱�BG���£dt�u�/SL��JTk�#���F++�gW6њn-�����JɟR�[���_����7��0�N��hke��O��(����c����`�
�d!/\��q���*G�N���,�ɶ����á{X�YBe(�en'�b�r�G�~�ص���O���8E]�J7o�i*�坙��rۈ-l6m���2��X��j�6h0��
]��ơ�ׯv�<�r�Ogn/�s��I�U�w]�8��.Gغ˥��κI;�YZk2�u}Ѐr>$�I)�r�q%̴�<�6�V��+7��,�7,�)�-qڨu�y8���P�ۖj�˄��4p�;8=}��)���P�4�Hι�JwV0]�N���8� i��I�	�����}/�Z__I�=^�S~�7�� �q��ܲk��[Z���?x�-��KVcOVko P��i��s?k�M�i-,������D��W��>���S�b�(i�?�`��x��@]�!pŪS������x��m�P�KNMMA��&�VƙW�d���;�qoV�46؍GT�Ȃ~����Qd1�yhZב��7��w�gW����v&I�����lG���.��$�B��/V�kN�5�<����T��}a̫��yM��S~�cG�u,6����7�B�qη${(���s�t�;�>w�����-J,�@%x�E�p4MSH��=Y~�8�]S�5`*-��2(s/YY����K�y�*3�[G��n0�:��d�0=#��ȒM�4�D;=�?��߷�ݍ
̟�aV/8���Ed�E�$e����1PdZQH�gE�z��x�{En�\{�陥F����h����R���Z��S@��f�����j
����fG[����#?��1B<���aǂ���Ҫqm�%��?�ini�}���4𛣃��A�!�%()@� ��_����:(�Ay��4�K�û�Hh����-�o��#Zyff�^�l��Y�8bÔ��o��؛��}T�D]e]��J��ѥ���+��4L8rz�	���ICWY���Z�Lidd�v���, ܤ�e�-����]���K�*31���U�[-��:d���#��inR�u�Kr�ʹ; esp��m'H�w$�M��.�U�n��%$�8=_�n�*��_����G�L��Q��_�j���v�p�|G���!��>D�x���G������W^�������tK$ @&�'��؝M�(�j��r�J���B��L����("ⶦ����|�{�S��w���_y惜��߾�A�!�|-���n�Z�xǔ��ŗ�;_���&!%��海��Z(���AX�t���!��O��,�����-�bŝq��_h��C�x-Н���PD,�b��zlU��l�Pp?NBH����=r ���V>�
�vO�Z�A3����Cb���o�Y�Ƶ�̅���-���x��h��)wc�4�ab5����K NA��r�����e<t�F�v��^E%bc�ΰ�I�<�}{�X�aH��d��Ǵ��@e��x�%s݁m��o���֓��2��6���Ol�L����[��z'��)|�Z'o,���:=�tAN%�ģ��qzR҃$��NcK��l�Q<��8���OI�c�4Z%��p����q45��Rt�vt(���ެ��Ȼ� �~x�5�G&����QN�`�qP&�5�
~ � ���3`�����H������z��?�P �;��Ͼ��pƭp���HͿ&Ѽ�ۂ������{F\���zG&|#�m�[�~�#���a����و�����7_%|��1���� �s,��2Ɋ�1��c�a��� �vAۢZ��~ �o��S[>��9��vT�z�?���W�f����~���Y��ny��b��D��t#<��@e�Ș��t��Ky����&����� f�~�^EY�D���G�\�[��I��*���2u��TwFF\��3_<�G[tG8;�D��U���
��wO u#!&���9�Y��`���� -�?���:,�n�4К�
��P��( ����3�	�џ�/�aBn�Zn8D'K�> ;P̑��Ǒ�륹��w���w�
uS��ux���
���:.���EI	E)EzP���V��nPI��K��[���r�`�������������|��C?zf朽�^�Yϳ�:{���5��s�����%���:W�r/��MZ�mѽzT\�]�4K{Q�8��5/��c0�ԗ(��sЫ/׵�r�fr�%v�F��b��{>��硷x$�o�IJ���V�X���t|� ~=�0l��L�D�p���zg3 ��*L�����>��pȂ�ٵ0����<]��	.��ƃ��}w#h(�����Ky"�M��&=\T�5��4��U|�f�f�E{>=m��7�I��.H�l~�ɯ�~�@y�����Oe���%���.���?h2�yTB��{��'��W�-H�O�J��/��� i���gR��3n����R�?~[��u�꠴ W�����L��J��̓��zо~�������{S�QF���$��}F,��1��k������8攗�}h&����3gk�rku��Ȫ���F�`��3������Z��G(K([{��hy)=�3:ﴇ�i6�'N������lv�]��*��ý�(m*��3�R�^��>@�`�ƀ�S"����B�	��+;���Ta��T3'��r]җP�WP'�����'�T�z>��T$�ƺ&U3Y�;&�G=,4��h�J��k��#�5����>�b[cES�4>h����]�!��O�>m��W�������y+�1�a"YD|�����!� �|� 8w^-���p:X���3�^��-�{�X�Q4E������P�B�%	dSe6� �����#�p��#}�M��B�l��m�R��
����%xR��ۃynFFF���s\~)��8�L$��Ohe|^��ڶ0y�V��N�x�;şq��8��WOO��NbA��D���/�HS��I����E���*�w��qa�&:{�P�^۸��tC�5�L�{I�D�r��׼�߳ �! :ͦ�L��QŲ\��Un1z��Mƣ##����Z��q�>'nG�8��y;�Q����ej]�˫�J������^X;�?�#}M�cwd�����p��L��pYy�UBLTT氂�<=Pmuז���'����:'���ӈ7��ޡ-�T�c� mC�i)�?����pG*��G��ӧ�L��"͆&7w���[���O�E��
��j'��a<�� h�0U|19��$�}�xS��.LL�D'C^��7���z���j
L���qu���|��
I�^�xR�=K7R����>������-O
90���m��i]į�m�=�g�MʊB����6��G���vww{I%�A+�4J��%�6ǧq�?�IING݀=@�9KJZ���8�­Rد_�X�}Rg'��:�PR�K[0�`��WL`�qʺ^8t��X�a�q��������{�3�É=��O�/��:�u�q��G��+'�q�=.���1��G:�W齫`t��_4N�HV6�:aET�����I�����j�L*^��V��ؖ:���ӏI�h0�g-f�~U��3`�}Ij5���;���]�%���*�,��VI���3��a�YeTU���S���cb2�ݨj�ǲtT"�Aj�V���ܘ�{����ƪ��(�T9J$�u&"bja8�42jq����?fM�D^��覜�%HGZ������}�K���I��5L<x}�V�å��.]�G�:��1(�W��Y��)<t��7�8�4��V.rVY-೘o��^�(�[3�^�;|�"1�錠J�]�RU6B��/p�r�A�_�c�{��3$�ʍ�I ���	�~�]�}	x|����4/�׷������΁|�k�?Qc�J���\�b����gG����ޫ)�����p�ذ3�%����qgF'#��0�$9��kd��>�O`�K��
�L��HrU#��^y�]��4����O���֖�����z�h�	XyY�ؘ[�du�NB�F���ɹ�*����[�z�˺�kLó�1���ڼ:8����*��i^s|�͔N���z@!����HXR����U���OXt�:^_��6k� �@,y�w����s��sk���^Y��2���j�N��\-�����n�Qt���C��kZkq�(>�?K�Z�n�jq�Kn����l��������?�9�^o�����%������9�p����%O��z1v�'�7�v���M�9������O.Cg����[�P�sa_)/�%���q��V���d�u��ͳt�����D`����O��k�PG��JJ[�V��)>J3���v�i�R=��l|tg�e��[�3Cpiι���'A����W�z�l�!{^�y�r��q`>����d�]8�39I���so�˯Usv�R�Z7]�d�[��2:��ߊ�|�	�h� ��'�3=�ȗjr��q����;f6'���Vƿ��W��!}E{�'��Bt[�׻�N�X����� 4��}u��$TI-�z�?�}:��w��ȁk#����a����T?���V:��4�j�b��.�24����'�	r��a0��)����X�J�g>����-M'\��6�Ȼ��|熿��΢�Q���f��#iY޿���-���X?�gs)����ép�B�j�)�u�n4b4Fq���kA�T��t���f+�%��U�of��`i̤���p�᪉ԗ�����ٖ�|���J|��m`�=}�x���+L���K�e���^����E��L^z8{�M5�.y:u��}�H:c�x���&I���ʜ֣P�w'3rRBy_��=a�\�t�;3l7��Iҩ�B�H6�*%)���A�!�I�o��u�w�V��h�[ux��������bTt�,IA�Oc����Y��;�//����?T���qW)Y~f�8f9$[�0�l����7 ��$,w�>Ǎ�f�D�Չ�l@�s�"UTU=U�E���M��{g�Lټ/����g�bG�)g-�~�?ռ�U��E$�++о�� U!��4vR�-D_Y*-
@�...D�i�w�sDۃ!+��u�C�;w����~�%	�ٍZ���
�;�z*"�fhl�;*	�7���ej��0/m�.���V�+WY�Ʒ1�:o���.$��*���aL#Ͼׂ2��ڻ����L���o��bc�lj�h��+Y�9��M�髃�I�F�o�y��{���|��"$&���{����1�φ�N��;��I�FM%�b�����-f�A1�H��ϻ؉�PڼQ��Ҵ��q�V��&���j����7�8���_�)/_�����iQ�XY!����Կ�*���Ƀ� q���6Z���3,��4�&v�����O��v���J��H6�y�`�:Wi��$s�:O���ާ]��c�TUCąDw��5�����>R���+�!�н�ݼtDRFfSY7'�-�Vn?�����î��A6O�M^�F�PɘW���M<@���[?���	�y?�L�l� �͓�2����]�1�o�Cw�Ň�՟��z��G����(E���>�ZrT��z	Ѭt��o$GG�-�����8����rYi�j��@'�i%�� !D.K��A9~U�3S3��7�n�n�[�z{�����K�J�n�=V�J,���ߍ�|oY��-7Q�J�x|L�c/5�(O�8���~.�0U�&7��E�2�*�<s���$���0�F>1�~M�Du%�	lC"*��	���Rv��ge�i;]��nt�)�C��	WX����
+{QOP
�v��-�$n��Y�S�*�^�k���9��s_7o����o��NsI��+|?�L����.����Y���Wn��W�D�r���-��~�?��2�~�W�q�?z���K0��Z�
�ʶ������c�Uo�QnB/����Z���}Np)��[��G�8j��x/��؞dO��nU �O�d���������z��w��\�� ���ͮVH�ؾ ��p~���m1�����<F��VTT��F*V�DO��d��[f�`�-z��<�t&+ѻ��v���0�cv���i���:WMuN-�	�>	�|PeEOP��ήT�d�pj��h����\}���1�NdБ8=�%��<��G(<�\{z��y��2�&1�U���X�W�r���	�z��Yz el�5� ���D�W}��(z��74��<Y����i�Q=�u>h�9��;MCI��t��C�R�b�X&�5)�[,�੹+RV��渦8o���q��7���U3�!���U����j��������|j��V ��HT�iZ�BU�a8�_��c�������p����;�ȼ��%���J���aEu�np��ޱ�-^0�r�^k�n���cq��SG77"n||�{�������;����S��S������*����&����{���-�f�:+Mg~d�:��S������(6X��r�YB�}t�Qo`���R͌o���F�0�<�xOoA�1�p�,�tI��s�0��w�ܱ��%�����[��M}�'���ͥ��'F����G�V� �@��۰3�c���KIS3�	3�/�꟤�	�²qX)�wם��W�C�smQ))^�qr������ ���x���g��&�}�&�c6�|H��(w�_�J\ow�F�(�z����k�(��.S�c�mu�p�^G���)#`	���o�&ѱa�U@��e�v��w[�zݞ��|E��m�W>��'���58X?`���|�����FnQ�U/��.~�f1�����\� ��F��bf����וj���`�i�Teg'W��K�J�����	p���5��g[>��Y@����Z�N쇯E� "��r�S���֧nn���Y�|��w�j�
���J�a ���o���U��������~���Ĕ2.Ϻ^Uaf�"n��;��",K��:?hEk|e�}�6�����I��w�˛�2U9��[����UX�T�0��hUY�U���~����%'<�82*���G���+<�O��CLM/�wBV���*�ף�p��y����b��Ć���A���y�iz���wI��սCz�T�P�74/X@���_�ȦԧO�h5��a�-�[*��X-�Q׾���i鲐�*��_�Rc��/UU��ہU���]ՇL�u���=<[O��Ii��P��A%i�`�ܖ�����p���2����脝���2K������tmjSU1�q͍����>y��f����l��3�[�.�q��GW/|`�K�~?����Տ��9�	.qa?���ٷ��Z���Jˠ���w�КG�wn��+i�vy���I�WT$@w�����R���pZt�ŧ�Q+�(Q]�.��c��)��u��V��u��ۓ�����\��eeY�J�ԣ)����o5W�%���O>�`G:�J�xg>�ŇxY�m����©������٦��d�]�k5�!TY�9kEHL�}����n�e����+�L3**}�Z�A`�҇r�<�^�p����U�$����}�;���;z*fTv�T���� /Tkn��-��9O�{��]�_pǴ��s�կ��U�&�i5� ۫n5bbQ�Fvq�_8���rU�t�,��~�^�L�#ү�pٿ�:CG�jc(���¬�~t�h>V�￟Ҍp!���p#EI���ښ�zn���1�
��y�OEU�8��&{q�D�4��M�����x����}��E����j)�k��wNH���AZ?-�֎����$µQ��Ȉnw�V�`uuU-I=����m�֞I��Ɠ�����j�(�����P�[Ɔ����q���nh�{{{}���2""�ߤ���%�j�3E�����wQ�wG��÷wJk��.�x����^�@~n��^���w��df��ee��M�܅���MQ�ΞE{���k�����9M^�<4*"�%���+��F9oL禥1y����sI��Z�i{'���v. $���}|x_@@���6�dg'#-Mʙ y�L��@%VU>�gf_��;��(��:.��zypp��D�����e���b
����_�@#��G��� e�?r��O��?�]goF'&�����#��SQ��x�jWz�{��f�|~<���R��ڄ_���ܜ����Z7Mw��дo�N�I�P+ҙX�)�=��m�9����{v߉�uGf'��죉������QuG�z������ǌ���i=h>*�3��һ�<����*�N>���jڟ��g��N�[X�ҳݸ�	�A�ŋ�;�i@�i@dOC9[��}{�͑C�/����)�i��u�7q�N�#�&��&Iv��B�9EEU�����B�Ӄn/� ����(��[<�I0'���f���������������C��1T�j^~0�B� --튃#9S��]`��9dZ�Q�U'f�'DF�M0�O����_`+8=_���4�_�d~�,%V���.B$u���-��ۯ��M���W2/��o����C�\�*)JlkcVV�*��gisم�$,����!�io�E���V����z�	c"��[�q�N�2�� �7���R���kk�c��e�CZ+$�cj=����h9�P��ust��Q�}آUe���X8u!P:��k����q�ޥ�ꀔV���7~]�ٹjk��gD��+��r��m����ܼ����>f�.}��^h�B����2@?�z#C�$�
Z��T�߿<�Z(��K��/@o�#�E�ҽ�����j����F�c��C!ڰ�ԍ0�"��|K}51-4�p��5#�9k�-/]���ch���v)��KNP��
�9}�d!��N��s���R�׃A?���t�0rX��G@5+�ܢ�:&q~o�iv�ꠤ9�^���.d���m���n� ����@+����/_�.�(e����-Cz`k�x�Z��	�w���}*�_+u�4Y�5{��_T�7T-.w�=Jy��T̙~���
0�D���mn«�疔��i܉��I2l��:/���:�O�*�W =q�N�#ݎ���Ғ��=����ٟ^p���l�r�ULսd�x.ݺ�P�`�-ˤ�/_RO�O�I��>`�lz�3��
듕�Sn᥆]�К��C�N��4��෧P#��I )CQ�衴agH)����z�]�@��0��36܈��
��Էz.]�!���S�=b�N��̲!�W�O�j�y+]��f�FoX�u�� ]���M�FA�N�����
��᡻�۷9�]a�3��Wi�ޖ~��o�+Au~�OZ���B��T�n9k5U�ɅS"��Ʃ[�BΪ0O�q�_�+;���:�N�b�r���~���T��{��jUUU��������I�ѱ16 ��1 N��W��һ/3^ ~��PO���UR3ȇHp�3�Z��������
�`F3e)�2���^5/�Q�V���C�S<
�l��>%�VD'�$�ynu���Ԅ0{��0���]UY9`S�JZ9����>��6��{��'�@G�q/��&Pp�\�-��'�74�TVV�Ң��F�{�]6
\P^���� �z�d0_v�5ֆJh����C���F��`����F/���ݝ�P�����";_����e�v�[��@az���s��жī,�C Z|���M�d���?�ߠYn�[S��"w~WXX���Lc��V;y����*���J�l�m�Pw6f���=
��J

���= ����w���(+))�,��0?9]�q�TQ=������|vv����E�<���L�$^_�qQ�}FB����v������w����W��^:#��(!�,F�����n\��[��t�?��=2���m�gn�	�[1�ݻ;�����f}�FXX�2T%����ۈ�o�*�k�L��_�:J�d�t0>;�3�Sե�-QM�-�k9%C���+g}S/�kЧ��K�9��ז.]��=�$\�zgN�뗰VV�t��7��żu���ro i��j��_�� ��q�O�����{v;wR���������>�w�^�Kûw LbaNlX��k�璄](��0v>߬�	)�
2��>|��-z:��.��^�DP{2�ל�yz6(����%Q�{r���ݼys��./���n$�}�1� ���qr��^+t��U���Â9d�z�q���n,�q"�ς���}�ǝ,��"�����|�)x<�(F����R�X|�����p�D��Q��1m�\����/m�w@��=�|�(�&v�� ��(���?Z�F�t���ՅS�l����
� �����@L�P�����b���n�(#��\�\�=��ϵ0�(/��KɅ+%��!�PX�㑜[J�	�%�---5���Lu�CL�p:
�N!3������;
51QQ�`�����㠋�ML�6��������o�V,E�r���5�T�?�:�2-++�	R�Ӯ���K_"m/�z��S�W��˝1�p�q8�XѰ��/����j��J�λ�[����R�j��x�(��|��L]G�c��I>��;�ћa�T�	�Vccc�a�w#K3ec� 2"k�lP
���钡g^v��|+�s�����f�1��`d|�����!��BF� |�?L ^`E�իVZ:��J��,�9�̴k��i)އ���j��#��I�&!��Dn�)4w�s��;G��h�|�C�R}(�>ڡ��#��e%�[=��Ҋ5<��ݑ�NUE�2@�G�.Z�l@Q�J��9���c���,=/�p �B�������8�}@'.,ۗ�TW`#�X�bc�Ԕ�ۄ����1��y�:�s�>��y�DX��T�Ք+�~we;����zt||�0*�35�����јQs������,��P'��N�r�x"���Tt��or���)�E���Å���.�tR%�xT)4}�;��]��J~���_K�<O�������J��E���sp*C@����[�^��^.��7�2|�_-�g��U���/�Ӵ�.�-/��-�ؙcz1_-r
�J~}�xh���Ү����Z�N�Mz��8 �%3 õ+��[�;
v^��i���ZZ�n�<�Gr.!����w���>v¡�ҥH�{��?��i�U��L�Id�~zδ�s�;�i��x�hzF�KF�]x�`1��q<\\$N����v�B�}��m���bb)�I��߿?9'��b���h΅�9�r�����4m�h4t�j"0
BR�p�P(��⣹t?�{��8��)�¿e�s�N/<$�䰫�7;W~-�&e����Ƶwt���̑z�Љ�y���6���i��BW8戠>�]=���@�Y�E|oc�F���/ �^��^�>y�k�3����Kkk!��+k� ;��5�,o�+��Ћ�;\�,1�+� �\:��p�spwv4�a�&��$��F��*����t}#C�s*br
r&c���(�gw�^�I\m<��4�Y�rK����:��o2>wIKO�FC��f�?Ho�HC(�@I.[�-
:���Z��R�B���U(��Ʉ���),\l��U�ɶQ�%�ٖ��hAj���R@-�'8�{;	;�fgf�x%O+h�G�_��xupl� ,~�V0P	���={���ag}��͛7� ]?|�z���0J55{�^�W��.���k�.���
�rw�O�����s� ���^6jt�R�E�r(M�
�G
�Z���;'����f�x�%�$�ݵ	° 2�����}k��d�67��޳��˃����30�S�T8=�VQ�~(å�
�@����3hJ�.F���U�����<r�Z\Qq������;7n�ON�5��p��z����������+��^�ʇ����Awp���@��!o�Q��:��w)o�x}�k�=	�2�ݐ`澷q5NN��zP�-/ﲀ�g���b&��"7�W[֝���E�#i���]�Xv�|�1`�����E�����@{2<�#K�ut������g��}]Z�]MBJH�RM- �tH��46��[mu��e�`]u���g;W������>	���>��\��{g������&Al{}�^�����Axy�v��{����=;����J��l*!{�ݵ�P��R1Z���A鱷1j��3YnBZ�S���Hq�w�1�������U�;���|⌬,�JcE<����f��CWWW��{�����'��lJ�v_o 7��ۣ �[ �'>v{� w�������)�B�m����%��p����)�|�m7��<�|o<uӳ�d�?b���P��˄RW���n���ږ�,��YP`��I����j����P:�.��c�6��!�A!p�ZY�wg`}�#8снM�����*�z���l!J�''#\;pYW2�	�!���`j"��pp��g287���H�҇Sb�
������'W��h0��c���&�����!wn������0X�`�2M8�pb)zq�������y$G�U��n�S�0ږHV��mmmm�[CU. �� ha�����>�QX�tm�n�$'7,�Cv���������##��q/w�3�9���`�h]u���ژ�i�Ǯ�˛�pw!E2��G���N��Kh�����ꈍ��.��p5�;`�-A&���җlQ������a 5nw�::n	R�}&$��>�`�(��B*��,�R�YK.%%e9UJ�s��ݽ9�!SW��1U�8�˟�\]ѯ4��C��u�L�����ăj?K�,#��|M���n��&W�~�,���[S�U�HJ*`��G���w���ed�ƺ�ks�)�M�y�t���)/5��0\|d$9<E,��F�JV���077�ô[+m��;���K�&ɉ� �8�L,�tj޵�?�[@gh�l�d&[�DЙ�S����x�K������XAi��]�D���g�!��w��llQ�-�
�Dj���W�o�8�n����o����372��_{��'�'S�/d�5εR���� @GW�*̔#���ԥ���⣢nB���̜K�izjiY�Z�璒���5�-߿|$g�333	\�&�z��I$AC�IE�@��c�b��]{jo�B;�<���9��L�H���Qa��RM�s���@3TA`��z���r����-Y��O.�%�[M���t�n�K��2Ԡ��Ρ*vZ�T5!���4?o���[[=�c�Џ�[7&���>����SH��flms
Pnmm�x���BoBm+����
x�ס�/�\�:riw}�0xn�K��o���hNmj�����]mJt��g��΀Y
d�{s��}�v��p:�:� ���68x��w��A:R+��@M�=!���_koT��U��fe�MJ1x�'2���zb$A�{zz�iC� S]��|���<� ӛ�f����O����F2��ׄS�]~�F���jH�o���Xҫ0=��3�!�&��,����p�>hu��p�
�b����7N��8����<�mC���	�2����a�қ�7�#��e'��]1�����H_�sb���
�\���C�z����4�8	�dn?������듣�9�0��z�ҕ)���,G����nZ����-��I1���"۲9K+���.6��<��"�$؄�O��?9 �"���3��o߲�$�n����7���~N@}Ǌz�l�.X�Op����F�i巖���4���! c�$3ܻR�s�p�FGG���Ы��v��j�p��9�h�

$E��a�xbfɐo��/��\0���Z1o��NZcb W�}N��r���ĊO��1cӵu�[@��J{���k��Ї��7c�
��H'��w	m���3_'A)_�n	�,6Y�Ďnq�ܰ���|R��x2��9�,��J��ģ���+��3濨�,s=X���#@4]/���Yn�][S�����c���_UW7�ǏWp����?�.j8O���W��Hy�O��ܞ��}q<D@��S?�`fb:���rRRh(� t���{7`a�d8�K.iQ�&|X���<�eP~"�!q�z�;��C�%��&&z�eo/���C}V������'G�p��]�@�R�ξ#��n@�1/{^�5鳘��&����a�)�	�c�r7�1�mS)�c�#--��$�4`���;�H:}ϭ?��K�1�������٨��4�H��Ųߙ�TJ�y�%���:d.�A�[ۇ�?#�"Sʫ�:�.5��1)��k+ �T�c�8uj�3����`.���ސlM:�&'���b�ܤ���4��8YRU����zN#�ux[LL�d{�r��Ȩ(��r` 	)��lL��M]�P׌
�Xx�}�34�k/#�;?7�D=}����� 0����3���-|���H��\1��jjj���������D�"(y�=y�Υ���C�vέ�|e�(�mH��mi9��y&"2R��<���f�)g�ŵH�%�],�D5%ᴀl+}�r�b��G�vR8 ����(w�9�������NAM��!���W~6}� 	�Q�bw��I��@ �P@�z��z���G��W(�ځm�66�9@��2黝��I$k=�M�q��;������CCנL�#S�ngu�nL���KH���A_X~
6�7�&M��Y�J��X�s�k��������!���}D�O�ѻ��ŵ���:��Xe���@n5Y�m�<�c�M8���1z�%A�]ˤ���[�ΖI�Y5���.Xd�I�W�S_��K@�tDܑ�]껕3j^ع:�z��`���͍o���g���АR��S(6��ŋ���.�\��ѬB�|��)P��ss����k`�6�П$L	������'A��ЩY��|�D�����S�1f��'��Skk�%xR��|��Y�vL��/����a�|;+��ٙF��o\.�,'|�;�]�VXB��J��8��oXi� ��j����[*���r�TT���$����Α��@d
�1��P2����<�t�L�P��=J�փ	�#3�|�� ^�-Jb�� pT���r ~�:<L8t身 ����H6��}%~r��K?'{��A�G�,�s r*�3�SD�H��ymY:A�0掎�'��fjA�����ٵ��>�_l��T��(=�f���k�iNR�����o�*,�/..�d�l�tT��B����|��U��V�qsr����䢨��ԍ�/tS��}����l#`�߁Y%%	�m�! Ͷ�����sj��ث��n %��M�s/���
_?/�>90aaeE�8
��>`zG��p6�t��1�����5�8^`��	�"�"N�*�V`�����i��5GG?�B���x�H��x�>%��2kܶ�X���h>���Ϊ�HR�.X=$6)�ս�ew�|2篵r23�;=��s���������J���Γ� ��8����n������EU�����!�����M�`���
^�k�%J��x�K�9n�q3xY�6'�xP &ܑ&�	\����A���t�+��!)*~�X�/�/��� �u!=\��Y�Lfk�5�H�#¨�>��7��8 �+n>����3� \�����Ic��*?D� ���9�&O/|�΅�_Ǌ�p��:�`o��5dc=��_�= rq3u�Y�4�Go��ɼ�*���A�A�3F'�Kz����h��yd+U[�U۵qn�Ǯ%�H�׆���S�a����X������S+lP�� R�Y���o [��D�TTn��
�~�ҙ]SC�@h���fm�<��Joo>2;�"��ʫ މ��|!r�QQsl��ZZ�8���9��($���/_�uϾ'��`i�KKz9�zpwm�M3�kU�ɺ������\eV�w�F:����������xر���x2j���&�lF�[qy���
�			%"h&G�q��I <�|��O�l�?�o�����(sX"����2]���u(i
iΛ_����$�.�Oج�N�rѫo��7wu=K>a���q�A��j��*+�٠���
�j]>?�mg� �i<����n�P��.�r���L�����g��I�vi
b��I��!���&&��� �uݛqٚ0Iy�n-v��p+/+�,�9�=���Dq)100<��W��
��� ����I=�x�ʂx�Iju�KO~�4�B�B\��#�R�C�b�}�f���� zT�F�+w��*��tm�HF�\ê�������Q{����-k�*�$�[��g޽��k7v���Q�^C1e�N@�_�Wn�ip5e<75��&|&�)��^n�\1���g�f�dH��_}�
6��(�0c0�b����ߎ�CI�"��{Fy�mt ЅfO�H���}���j�-'�vj$y������mt�y�֭D�]����}j��;@9~���J<���
�ӠmF�,,- 2'b��7���T�y��.�����^N��8���ps[��v��ū<�����E�N�+���	�f9�[!n���8��K�AW
9,Q	R/�v� ��*))��׫��~���Cp54��YӋ�" �~r��G�9�D;:.�M'�~��{hq�~�7b����t=4_�>���9�p�7'�&vGb�
� �KI�MَyD���t�/@;=1A?Ή<���}�BA3QI���fE���,�h�RVns{b�����a"��^r���L�1%�99�~wո�����(��������(��:ill�dedʂF�xս�EM܊�w��k{�,'+^�ح������1}��ť��!���wc����u 4��C��A�
��Ǩҥ�%]]ѕ��[_ۑ����� Hۺ��d�1u(!d��H�	T��K#kS�=����ϝ�@xW��ى*�����#���J�$;�-�b��.1ec�|v��w�7ơ���������u���?v�N89A�n����7h��w� �s N�X���^(�5ve]�ua�ggT}fL�9;?�*����$��&~ � c�v��O�"Ê&����� e.�g�@.������˗d�~zp�l��y�.�Ş�*���+��n4�9v�P@�?P� �+��p/�h�*�B�c,�T<Q��j��C�R
X.�MR9 ����'���u;��)�54���霔������|�]��K�3��BD��K77!��9"?W&=L���^�?$�n:���O=�i�F+�:�@C���b�|�H��o��P��zlS�o��ɼN�o�N&0aO@�Պt.���1�ќ�Yg�gffn5ċz�!�k�;
tj#p}����n�ڪ���1v�In=�+?�=!�L�4r��ֶ�k���٤�?^���bߡO���1!���LAM��&���b� ��s�c�gr�H�ڨ�&\�(�Sa����DD��/Y�;cFQZ<c�ׯ����ڨ��+[=m ���ke3_!�����z���
4Z�8��.�N��0x�I* �Ez��s��v�1k��T���"���ВJ��h͒�g���联.h���8��B���Y�y�k)����Ǵ�Ra�Tۨ��}7�LT����	���aʃ&��@'����C���W"��a��A���!��Z< �D�H�S�R*�� � daRx1���[,�a��^�|�B�Ց�ϥ���@uAt~6�"����ʏzzzN=݀U��p�p��+B*g߁DM�n�:xmu�)�t�R��C��bnnn"B2����Tu��d]��I�Gg��2�Bw_O ��E�E�/Z���:����h b������`N���(��c�.h��"���t���P����s�X�4WE=	r��l˹�~��\����4h�{m�K��;pA��m�$���*��X>��Z*�5�S��@^$hU�d�2�Ł��Y1�ߋ����fʍ��ZZ�	ߜ%���?Y�nd�}嬒��vBD6T�ز��r���v,j5^�:�Y>I#b��yM����Ŵ���Z� ��������Z|����K�Ƨ&���C��kjj��CS[Q11�[�@�:Vh����ܚ�ZD�E]���7ۦ���/���s9v=��� ���}(�k9��]�Aw�0���+�@Ȼv5���^!%�q^���^���\�a�8����x�dT��Y@��_g���EzĠ��'�1�Z��+��E.��d��-�ݽ,���5�?p�X��f
����y�w�qд�������g�g�����<�����\raee���E	�Ё����!�U7<Ydj��3ƹ?���v!z��/�+��X0�Ty���ar�&@�Ƣ��r����Y��^;7����"/\��x"J&OyɅ�zc�sДX��l+A���/�`ýd��&nv�O
��7)(����=�VL���VX�s�G�utH`J
�>�As5���c�O��>V��|$$�	p?$��� +�F��,D��ʪ�
p7�\�Pze����\$woO���1���BCgGǷ ���bA�.����"N�䶤{'�x�ChG�j*��s$�B��ӐbAJ�P���r�:@�,G�45���EzNv��Kkj�p�,��,��8i !�֘A�@�μ������&"~vg�t� ��.�����j�����-Y��}�?�����Q�����2\K�i�v�N͗_t}���~ ����p390 WE/����\��&�K5���⢢Fm�Y�_ZY��`H񾦃�B������?�1>N4��E}++{T������w�h�L����5�"z�p�M�ְ���]>0}͡�"�###�௒�@�r@u�mll���^^/"�?��R�����454bǶ����ը�yB%���Bm��T��Ui������߇@� ���jH'U�acww�H��W���)A�F����a��[���p�j�ҙ�\:/S��.���o�I����S�S�b'��o|����O�������N�� �����{�.�xH^���E�;� �UR�_ߐɌ x�X￤ȕ�����$+2e����������t �8�	�8[]�D�NNN醨;fО�ɠi��S#�ʕ�_#�����:X;�Z��1<Ls|xt�9��n5uxjVUM�?V,�im��a?��->V�lBKvV�y�����K.���Zؽ��#9Jx/ ���~vs���a?8�\J/�O���X��OO7�e��K�����c���н3�>���=o�V��ca_�H�INA��|M���y��5FƧ�R@@����֦��%�8��෱���䚦���;{{�'�HSD����p��ēu���5&&$o�/_�:��=ӣ� ��ɕd�r�-E��!^S�U�8 �<>� ��ecz�S�9%Ŧc�������|���=��
gX��u �����)-�^� �{�����㻠]X��l�k�̟�T}��V�����,�(~�ǔ�����E�Ra�Ф��B�ت�Q|<��nVST���qjm����;x�0�Gs��ƞ�MWYMA4@��Y�Ɓ�� aG��<���F�q��nF�g�w0�$�d��Bs棗ec�$����E99߁�̔�tČ]�BL�� �\�]����:�����Z�4s�.(/J`H�@��	!�����������B��Ie�MU�67�_d{Pa�%����wwwww� ����=���%���f����ݪT�h^���9��~��~dl,Bn�����'�&�5,lf����n-� `K##!�|�"��6q@��bcG z�DU4����, ��o/�g+������P|�gO��wD�55O���W^ǁiA�Ύt�x�j*G�ְ��rg����^_t"L�$����@)n^��vϿC���Wµ��������������!N����=b�@7��\�M%ees�6{�1�h��@ȋ� llL"N�R4,ȟ,6�:�-A^w@�F)�x,LO׮�� �y�:�wB%TY99]�h�����v�ԸjY$43euUw꾈����U��%�"���5�9��TlfsTYz��	gJ����x�KQ�:.�+P�}\�1�Z����������
����|^"P���p��y��目���ܟ_z&ΧK�z�@��|^�_H��͹���9��~vFoo�y�=�&�%�/Y?Ujk+*z�𹜏fHj׃,�u"���Ҫ�8m��}���Ncjj�}qQ���Ȏ���SNiuE'B`�m�QDaHVVW
�&\Nn���S��0VQg'�7�D�~�@��%�euu	���mB#xyu�oqK�����ϊhhh�]]� ɍ/ZycF�BAA	�~zy���$zxxH�-�a`����
��Z���t��]?��a���ass���1�p�@���� J]6l&������JL00�OW���i0������=���0��H � �\�̂ȩܕ�r?����fA+w���@p ����
!�7��������{ ��������$ۆ�?/����� M��:���K5
�5cQn�\U]k)�P5�����.)!
�-��$�$XQ�%5�c���Hq�P2%h4{_��uW��ٖ/, <���/�Wܠ*̔!Z�
h\�6�0���Ly� }����6Ѹ�J���?x�y�%��L!��p�O3?+%-(�{�F�Ui�T�����E��m�8D#�"u���M�`�l��ki�z���L.�:2=8�7���¶��U����ą4��E�r���%�N���[`��u���ޙ���ɂri��u��LN}p���C�kG�-��\�������EF�|�Ӹ��,5]��H�!I�!���q}���R�j��Q<RK]��pA��N@�R�, ��0�4F�i�ο���|ג'��4ԩJu~=�7 n^���I�(@������X%��I�����7Krd�I\���W<��5'�l��ċ+�hKl��JS2Uw�����E��L@\�^6��Yg%ld�9HR̎e�ߎr�㎨or�hqqzZ�{v������������Q����v��NӸ�x���e����Z���T��T�=�����j$4�A*Խ�4�
92B'��Iz'�?���?2�� �8�4ٙ�i�� C�;Iz#.����٥��T]��R����4����6��w��m�0s/�y�NN�[�M�S��,#e�H��*Efgk��4h�FR�8��ɖSˡJI�-15'�xO}= 3�Σy��`za��� �NR9�ZwY���w�n�Q@@���!ֱ���&�+.��/	�~o��յk�c�������u�=��/�5	e�$��ݝ����m� ��U�c���}�������O?-����ޜ^ֵ��uqq|���+�9)+fԣj�7<Gnb�P!�Ɉ��R�0�7A�^#�}8���WG2�h)j.ob�>Ɍ��#�hM�vaW3�@(�)���Xi�V���vW'#����G�7PUP?�I�	yum��K+80	LI�v��w=�Tش�ʇ�3I��T�>�❕~�Ae�Qu�CC��~��P���*srx��{�(�D?C����Κ^�>}Lẖ�%[k���B
����J��&:)5':�Cə�4Lv-	��]/ ڧ������RewEB	5Z��z.�1@]��|!c�A�W�Gh���$đOyhꖚ�LrC�1Q#�E��{~��Q�	c	CL̪1x	�۲��2��_��|�s�I��曽��G!��!��%e%�/]�=�gF�%0�'C���^$���c_����3��l�����Ұ\^I�|9w��0�-IK�)ف�(&Z�O#��P^(��:8���.=���v�7A����IF<���`N�F��^���t���h]7�9ð�q�i������䊡�n�����ƒ�� Z1o�W=V\t�58���� �A�>��(J�+����,����SN�&I:�3u��;��/
��%����a������\]��jfJ�X�Ð��!)�x`˦�f&��)�bfI��YsEg��-�<� H�^
1^��c����Rha�ޝ�+o�.瞭��2�8 21С���T�ǫ 1�b �G�=�B�� 
tc5�%ҷ1�~�hl�����-&�8x؈[�C1e� q]��:���D�ي��y�(
�㎈޴���2�|:ev&�
�<)'P�BT=T(����ߦ���?�(A���=#�1�~l�)�X
d��"2(�3�e�c��%��ҡ��x�~���a�StD�'�f;��3����ڶL�~�BcݎhP^Q�Y���J�C8B$V�
���\Q&ݫ�_��?"��kw��(|\����C�9KK��؁K���gq��z_}
���
�;�8�~�	'�FGh�?�X!3�6�CT$����a`;����l�/��+�?�p:Zn�zn����V�׳Mi'.�5\./Dּ��������N����`fɡ̏^�Y!a����,a��lZbf��S¨)�y[.g3 ��C�@F���X���6:�D��SG�fqx�r��@)��~G�Z�b��#���dc{�Z7��KB�+姧��
s-�~�q�m"ΪY>���W�J-7�"�߱����P�B�Gd�1��V���v~�K�aAʌ��������d�yg��������Ì
���'|]P����0-m���שݾ}
:7c�u�sVOs���kL^�.�؝�4��߇���<(1�Gs���b%�0�����f�?�\�~���:��\h�ꞇ7)`C�V���sY���;MqԀ)�ϣu�N�X����]I�f�������m��<!���tl@�hȷP������Ŕ��p���_�X��Ak䝹��<AO��NQ�ym9'ly����σ�������I����b�����"ib��De�[NO�Ė��V*��Q�j����*޿�alٖ���5���3R� ��fz+1�$k�a3��Ȭ'l\f��AV���E�t�iƟ���׿X=؄P�0k�2�?�T�tԎ�?l���b�&5Mh�YQ�@l��Hd/�1TuOERN�\�(���ע��Εh���ֻ4>��Q+m�]�c+�`��y窤�K(��20~���0�.�Q�#EJ^�8g�=6l
���Pӈ}t�ݹ�����f���iص�Yi׏�g~~d2�4�%������k�ZYSQF�l����T>�9�5NC_5�^Oeb���t��_ݙ�/p�i$���Pد�å��6�{���ћ��/.�f�1�]���Q
C
c�YՍ���B�``W ƊZ6�9��au��>S!�4�"]�LN\N��O��n2� ,�Q��y?P�m���)<�k>��^Oi�;���A�RB`FY
pkɿ>՟����?qi�C��a;�v|}b��yz�j���֥�5�����n�F�r�ܑ��<�] �&�Eմ��@/�F���f�!���j�������l)-�$�y�?*�Y�G)p8��_�Qx1��g����,΄��������gDP
�8e'�ƅ�mV�8��q�Pߥ��'�ұ�ɛ��}c!8s Z�Z�v?�,I;t�`/�a�,�9�V�#�䈓�����=�]ҍ�W�"E�S�w��T����K2����:K
,��I.�u��b�N>���������B��o��ǁO��d�㔿�f
��˫�z�ʩ���s���/N�,���4E#L� .	�DY^E��QR��cak�����f'o�P����i�u����K����=��r�eV���ul=�?VS��ğa7�t�ꎹk6�I�i�� 8_C��av����}2�uQWW��-��x2�y����Y�9�TQ��\z��B��ç��]F��tdFƭ)�ؓ��Ú������_�^TW��U- �_�R@x1���'WZԢ(a
Y�,��1@Q��Ӫ4 �&	Dﺮ�� ҊNT�	v�p}B�v$�n����)��~󍽠�^�����?g@��F�^�{��^i��������iт�JH��l�P�
e+C�����[�"aV��j1'�z��
H���8�	)��ۢ&]>�"wfi�&(;��Tr*^H	�lY%;�[X/SNS_	��el,���R8�sPjh�uyo��y���Y$���������L�40Brp��M5��Tx��A�.83ɇ|�/
h���%¢dO������B��������S6�]��!�S�I"�F�t(�fQ�E�[c@g�Gw<Z#r�3#S3d
�)ƫ�vU��i����^�~�����ęi�t�?�X�{C0x�b2�&K�F����P-����4��{{ڪ�?;C��}|	�(�3�t`�&�Dr�~���0�a��A2y�70�?����HZ�X���t�Ë4�ӚH )9r�(.���O��S�A���'�-� ��X]��Ur�%c;�1�qH�HY�G�lT|h�/sgN�:]o�� �ɀ�)Q��B�����hl�B��(���0�
[Y2��1�� T-�|�(6??G��8��iǝ%I��ݞ8�.�����:)����<��G��el���]�4�l펇�� �W`�"�Z��KA~n[{3qJ]�#�y�8�d�@?���C�:���m�K�(Cc)b��g
$*�y��<�}I4~)@0��9�u�<!K/��ͻ��%�$O@�5�(��5��P�P9@} ��P	�h��,zwzM����T���
Sq����s���"A�����m*Ol��\Ԝ�,'��	? ��M��H3� �I9���ҹkJ�!Ma:�-���1���%����/@�~	�M����>K��)2�������*� �`'\8@��G�.��3���V"8B8RI (�J�˷	�����	܉�J��g��i&0:q���0�+籁qR�ޑ'����:U�ySS�A�瓄�u�%�?��7�}�Y���i>�X1�+-��_�)��,!�%��bw�Tר�c�G��W����L�(s^���i	�˱l������0��?^�Ώ�R�HJ?e$�ࠤ�Q��h�	*�ߎ/�UiH�M�osS��fc�h۷C�h9�P�a{@?A~3�fv�����m��ȸ@"65_'ǡĲr�q�g���	 � 9 Kl��� ���͋������0z���k�; ;Y��w
��)t����'�L�-�g�'Ce��'d?@����tU��O4jG�0�x��s�Ί�.��K���)�K�&��ͬ�	��4�)<P�n
��q�d�D��#+��sfWi=:��-j�0D�q�/���# I�
���� �ͳ
G=�Lcn�6��Q�!��K��Y~s���D*B_�act��7�r���t!bMay�K7h��� ^��T��ה6�g���= �I�a����+��X�IhU`��.��Ю9Z�����L�' |����A��l	AA� �k��u��N��ɀ?�,�R<썈����[����3D�2+Q���7�wS4v�Q`��{R鲞�Y�h ��.����}�}�  ���F���|&}�B6���V�X4r��R �\�6�[G�����: ���&���}�)�8��>���4G�#_�s�B�[U��`-���K IJ.�B�՞ck/B�'���|H�rpU���,��\�0|е�5H�TJtȁL�C��7�/�ƪ0dI0��wy��"��$�2�(b]�0c��`E�Ǣ��������>��Fm
 lu��@�P��b�f*
����7�`"!�dy�^;��|�1 q{��5f cjrv��(Gk9,��=nm=z���
�!4q�(���s"��$�&;.�X<z�p�Ӥe��
�Zv�^gd�u0>v�������8�2 ,u�?�(� ���t	�΋ [X++>��wa O��p@�*�ƉG!��N���+�\oH�'!�˧��S�W\^1�%��e�8�a[������ɨ#PA xp\z~���3�(m�C<�޹�FCBq.��ύ];��I�wD%�ZQ= �%��[gLP�}W�~�
�� �
8����t,T;�w���� �|vCt�*�GfxT�j��{J'N�_�A��nNC�R=��_��4l9�i�~V��۱�Q�����mS�I�`l�ܯ�W8du��r���UjK�7rh���1��(<�-�A�U��R)F����A`�bE*���Sָ��ȴa76o�������<ܔ�\��'�����4UJhk��4�����ɲ�ݗ�������F	����;�1[D��J���%�R�q�$m�l�:QR1`!����������dI�%;�5|L���uo�Z
N���~� $�+13'�_�*��6-D�p [R�k����>����&=}m����G{C���E�U�m����|`��)��BU���\{�.�{��-��A����T$&��-�
�7V���ܼ��9KB������I=U�c�,����(��2�%���ō�"�Dhn.��x������Q@`��O��~��o8��O~d�2�3C�Z	��Y�������L�Ƞ���?_����rG�ԥ}�L��Nk&[_���,�(j�%�p�w��P���P�z��i-��1a���)� g�k;����"Y��MW�A��|OfJ)��Ȼ7|E�+�.���A����ncqm|tN����h[�c�)~�0,T5L��E#fi��|,�uUL��,��5��J�^wE<7��EHF�k�õ�����ML2lL��-{G���g��<
���V�R��C�����bє�ﺪ�.��'>�/V͒�|�~��Dh!,�LI2Ť�o�k޴ =p: I\���1������˷��Z��H�<<�&���67�[���g�W���2P)�R�ts�Lr{|6d�7�/N��\��=5�V��X�n��L��<#����|���(Tt��j��8�?��4ZZKd�.����;-���N��ʳ�!Pk?�<��P�������6��#_�W� 3�	��C���UM:K��b�~����1ݲ4����ke��UX�����W9��Y�ߘ��:q���{�������x��a��wb�5}�����J484���E�X���MQӷ��AG?a�M��	��F���!�OG�s�����c_G'��Ɔ��12��G�/V[�'q��5&b�>v��O.lZ+e��HIR��W���Y!`�bp�鬜���9��Y�S����"�u/X���X^�7rsi�ǟ+*a]��<�j9�gtǑ��o�X������73��G����ɉ8�������mc���Z;d�2,�W��B�8	ba�, ?�O�!�O��X�5�5�_��R\oะ2�����K&�y\�3����O/j���^�}eK�^�l?v�}�����c���Ƴ}.���NI�S������:�Z/S����v?��p��|�M��kRt}:p�o��:lao��@�cPxcy�L���&g��;���Y<�/��">�5}t�N�J5��JH&.�;7�\�7��7�u� �l�<7)���J�� x�2���:���$[C����`��k��Սs���� ����E>o:��4��I�P4�̣�S�6�F�a�K� ���g��_��F,^r*e)����Y��t��?�}tɊ���b��i&:m �]�����"������m<8�~q�!�B�e6�@���m;�J�v�E�̫h�Xz��N�16�]2���,�n�;{h����r0�G�	 B�u�z��lX�1�Hh�PM9�q����*x���#��-��#���y���j4�4�΅�|��NC	�҉.���Y���&�nV'x�Z(q�p���L�ݺ�v7�u|g��46���*�%\]:���̾}k���+�\U���5��A텠�N4�!�b�������-���V�F�N��?�7�Iy��*\*�e��E�u�(������n�D���j����t�t�ۅk��ۤg��\�D�҂��[�1��[`�������Ą���+#�Üo��m�M�?��wz����qd������V+To|���~�� m�0�K�ВO�^b3���ߘ.*���X�:��)f��p�÷a��7�=eX���%�w)�i�x/�*OhL!�j���u�U���fæ�1F��-�h����T\�|Z��x�T�e�����&�aV��SV���4H���b|βw�BGl5V��ҍe���A�-A^Bb=��tq^'e��-�H����x��@,���j����]��FM0����/�ڮ��7:���/�}�1j,��+u��ݶO�+;�f˚Pʩ��ld�O>q�k~��s헳ퟵ��)}��иTH����Z�u��|gJ�z�P��k����ӫ�0�C>�c(V0A�#B��G��H�cRi7Y�U�Y�����]Uњ_ֿșUm�?y鼾�q��U:��d%�����Ҧ����b7�����*}��a��~��2�A����f,=���*�$��ӓ4���Y���t��٢L��
�\,0a~OSE�"t&R_��A�盹h��޺r>����֔՜��햩���V��
x���bO2�$B$ѵ�E�-T��E�:�=��:���?G�"e�̸�z��,�LWB!F�UO�]�9j�쌱�Z�8�u�(3xe��Ң���'���SR�p�������2�%v[��e��b�4��p�"q�b�9lx��D-D^T��J�	m����rG�����J5��z�ɩ��������z�]��o]F=*,X�z����Y�\�b��w��:$���!�ĺ��	�j�.��R��x���҆_��5h�<��F���W�{�.��#��Pe��k�PUZS!M�g�4�H|�v���l����}���yt�@���)��R�h�7�ɒ@�	�ԗ�e��������+�`$'?�	��V�vw��Z|�������t��
w��%�,=[��?R�#�9����92s��Ě�!w��w
H5�����uV�
{���;�<���M�fҡO�[�)�1R��̹]@y��a��\�:����yO��v�l�Z�\�Z%W�K_�1z=AU���szD��(Ġ�e�=}�2����VDK*�dNp�U���A�3���Ǔ����sۓ3z�j_]*t�Q�]{��qS��ՂD�	Yv[��m�	"�v~e��q����7�5p�o��t���C�vwg0�Ò����<��uH������Jl��j�e�=�����xY���G\?9��Ȩ��͈/�7��g傟�� ��n��*z���X�`mS]cS�'J�l�:OB��=�I��=�'�����"�/���L��D�?s����F2�Z�_|k��.�<<r9�<������.>e�S��X�}�DC�g˛/��e ����}�	KW�WU��BM̧��+�P��޴�Φ���7	���i<���܄,��������������cH8TLJ� z�{B�~�}J���>o���<���<�d��	mJ��)�,�� �~ڤ�]��O�Z�i��Ά.�
����	{���D�z�yX=�bQ?���o�5}��[�y���U��v|��LK�$rC�c�dI�G"�t�"N[,Ms_�0�E/04{�]��k������5ݦ�el̆��2��T�m��O1mGk����5KHmbh��܀hO�B]���?<c	4�.�嗜Ϝ�/)T��D�hX�K�r���OԶaX�x�(�'�L�{ĉ3�E���u�n� �����0�I����D��WB�z	�
��*�"a:�vOp��x!v����R�!_c�C�X;�v�DƩ�r��l�H���udu�()�����Z�>2�J���Yľ�B?���?^ڂ�\��P�x�TQ���*���I��
�?6-�^n��o�[]�}/r%���/�g�fwU�i�4_hg}��i�T��yk;����u3�o~��n���»�Q�M��/����1MV�}�a�<�eO�%�B9�/L�A'���%zsAM���?��{�.�*b�I����wWpO�#Y�h��<z��W#FPf�Iu��[��8z}�*��q�����ƶ+�j��cH��a�<�7h��BN.���d�w-�L��^;;Yz>���Lfи����L���&���	5>�;~,�-_��ಽ��=�aD�pOp��4��כۋ�����\��c噘�*=�'0��z�2�z�7�gWnM�v~�.�eצk$L�~�u�,'5J<���NzJ��l��E�9>��*�3�C[^И�������ʿͤ���:���M���.{R4x�zǄ4ѭ��|��^�"]A� ���,l�	+�?��'��P&Gl�A������v��`��3"��j��C�c���K��2��͝�~,/#I_�����J���ihjV�\S�,��*�{�HD�#k����Ϋ��j~ �)ڜp�/KK����wFd*J|�R�`ٹ��-���}\	�;rrL�{�L�Z�|mD\�M��=�Цc)Go�t�5G#��t�>��>��!���&�F:$��ԙ�e�W�HR�a���v��m�1���N���!o;	5�p�fc����F�1�����-zjڳ�Yv��>HG焞�K|�����"�쫊ܷ$����b2�(���F�B�d��B2�	�K�U4ݝ��8Y+��8U��K��=���� ���V��~���	��p����]����@gz:V�B�/���@�2��ؙI�f��K/Q15jد�~ov��$j��ͫ߰o����?(P�K�}�2���UG�RdG�8�N����o!�<��%���r��fӪ�2���y���4j��|�˵��`��( v����������1C��>8�%��7����S�� ��]h>�l���-��\�Y�;d�''U���m4%sŔ��:Q��ty�k
�N��ӓ��q���m�@�gN�
SDk�D�7����^3�-(2�,��������_R��c�8,��K-��|�^@��쿕�Mj&&RMYcq�D`}���2�vb0��&��H�[���j�n���K�0�rv\wwH)�e��!ۈ�j��M:Mv'kkt'C#�����������#��e�w&PD�q
�g�G����E�s�4l�������ɝh&�]��P�xi����&�y�j��|�U� d�>���4���^��L����c0���ȇ��c�_�����d�����2�p=Pdgl�S�������j���Q�*�R�l]H���������<B)�$���i4�@/��O2��d�K}�{ψ� Z}��$�?�ҔZ&�%;�K�<^Ȭॉ7����>1Y��u5����S�$%�����b0��M�[�Ӧ���/|<$�a�ԛ!R ���N��MC����9v "�n������p�5��)�ܗEj��J�%�f��h|��1i�'��ikR��i�U�����=����l��[c"�`�oK~�^�N1��
X�p7ׅ��֓>%22AĳM��U������jJ�,���R}5���H���������3�[$���`�f�_�d@^�ܛ?(b�1.�>tu�G>�'�����=˜�� $-
Pd�.�]�M�c*���K/� ɋ�1u�ߩ�`�ŕ�γ\�]S��:�h�q�%�Ӵ��t����=a�d�q��y���d��<��"��W���)�#���
q�{���S��{r����A@����;�8W���|��B�����I���c���Ft��3C
!ل)��҃1�����/�m�nt�:��nF$*��������D`�͓�`��Nd�P�T�5]��I1�^v~��3b2�{�}HN߾W�[)��QY[���z��3�_Y��YE���wxk|-J�KH��AҦ�
gG��5Ă�aT��k��53���Zl_����q�XT)�s�R�F�7�r[��@1k�A��>�y�L�Vڮ��y<wn��'�$�M���:5��,`��gݫ�Ĝ�#����j2(�j1C,�n~�]]S��"�W<���=���܍O�C��Y2�A� ��ә��W;6�����̬�f/Y����� q���C,Ӳ�-�cM_�f���X�TO��t����'LE�4��l��^���+�v'H����}˱q��<�\�@�xaOO����y��t8�$/8�X�$,
-z��N�����0Tg���d�8'�ӱb�L6zoN[
0I ��N����s^�Q�C�-�����!WT�˧���O_ʞ��t7G"�p�%!���fj6�2�;�k��1�U#�=V�hk$R�����.��.�_��l�w�gQ�%��d���;���_&C(�_�L�3��#'6�`Ll�d<<<?NV㛑��o�Y�C'�@q�*v�k-;��|�����/w��&(�j&�4�mj��ֽ�;��kW�t@d�T�nF����0�%�
�$*��,���c:���Q��~���0+B' ��&��AB��1X�	�e1%�X����YT��!��ӧ��������%vS><�ۍ����ĭ�����H�qo�� ����r�:�����E%n��=��]��i���#���Ҫ�;��p��W�ZX�+H�{Nƃ�pW��tVY�]�O���A�]nDn���J�n�*S�ԹKA�9�Q��%�v�N�乼���]i��e0�����;�D���o���1�䬓X#���"�����
��Q5����VW�8��_�JXS�wWg��0���.Z�=l2��ѹ��o�Y��7h������z��o�v��D6�Q��rpe�w�$���M�5g������ԓ��W9�}��B?����<9!�f	&80j"�����M��v�xr�K�h�{yݛ��-����
��2�g�?I@�'�Fc�]��٢TBQ4��QI���wVY�$N��ħL���s�&Ҕ<)5�Cr����R4�
q�$�6��jp���8:�̷f����ٸ
\˙@]��T
0�2M�5dp��=�z_��<>����H�(�w#��q��^�?�4RY>�yE�<l��Of�D��ː��"���-�����U�k,d}DV�#�9���ˆah4���'>:鷺]�8��1�a�?/	/�]��"ND"�&T��m]����p=�syh+
,�����]v>q��`%z0\�S��.=���)�F1$��p}��[wy0CAs�!�rvo�F�[����7�&pc��U��.���!c�-M�������̙>�L\4�6�V'�|���bN���^��ObR�=8��,g�uK�y	�nzFʔ�qs3��d�?�G��P'�f�|V,�������VYB�oI��2?c.ZB42~`����M#Q�����e��0q�:�������w?��ow�g:؜��#�qd�Sj��-]*Cꈫ�aۆ[|&���s��4��7xsW<��&���+M�Ia/m<Xu����/� �[�_�Ԙ��@LU��l�/CN�Ĩo�B�����'��ߋ��O��P }�Wg�]h����9�鱴>Z>R�U�Ȉ�q;�{���/�p�rY3�}$�]f2v�GX��M���|��e(�i��x�5mr�x(���o��#'�mF��H�?H���D�'b/���Y�M��!T��[;��ë%������^^��co�cZ��M1CG�L��3a�ZA8{!E�ÎhФO��5|�d%37j[����4g��ۮ<(�a\��E�z�g��Q��<�g�[TRF���e\�t��YZĲ�}�>\��|c���z�����>���@:�-s=��WQ(}�T�wM��z�2}��1�I~�e�,?⠧�B��Af�X f��z��9)9x��S�n{�3#LX[5k���d��|;J��O���PK-�ݷkz����UY�?��.$�[�싶x���4��S�S>�o�3�4*�:����y���T#���PFrv^���"�m!j�z�w�H���!o=�bV@�l���<�����k�'��64ܜ+0��gfC}�n����&H�~�5Cb�켧%Hl��L�!&�ǘ�us{{^^���*���P�� R�L�1˖R��"�k�,�����1�=��?ELF����g��b��*� o��?L`��������Q�}^��I�Y��z��'�22ѤPՈjCcmSK���1dC#���KDȯ�	n`��e��A�t7�Z�hh����+������\�����O�P)Z���rF�>0n��g��&/±);�J�R��9''���y�t_��wB��wOd��y6(��>@��"�[Q����3�6d�ĸ&hW{6�A��	5��c��im�PV�T"'G����k�y�����(>�<��e�&���n�췷A)G?Ցse�������?>&�\R��(��[J>~�ʚNDl����ż�{�~�2��Q���$-r��Z�uv@[Q�Q�#}��v��~4���~�/"~ߢ��=)	�S�=��������l�]^#.w�&��7+]�~�5�]���$(�����cQ\�#���j��kcƼ���P�Hy�bU��l%%%-�� �v���8wm��;�����bbE�+6�j��ճ.e|2���i�Dͦ�<-)-�UϳhC�����~3>�/!������#�q��p6�GN� �\l��SL� �J���۱
�����뽵���6�n�t~:��'n8�Z]����R�/���;���釼BI*��7��&�1T�k*�o�����+$�s�djm8vX���@C�����Y�
��~D�J�<0>(�#C7�)B:%�@��1���s��<;Gv'��@,}���Q$��*��<(>�2n䛅*��@C����[?��h����5>w�\0���}~�ozl�i'�Rk7q 󲹄^�3�c���+��yzBL����� xJ0>�(�ن90�m܈��5�x2vV!㉃��	�*�YR���佂��d�	-�z�3�?HAې�� ����=ڔ�����(O�`|~�Kbd�����F�	dg�.b��(	�G<xXӭ�^�S���<���_uM�O�� �R��N�N�}��djs�xĈ;�1�3;�/Ԥ�YN�a�cIl��:ބ)�?;�x۝wֲ׸F#3��\S�������ٳ�l�MA��VL]$���ك]�B��]���8d��+��HyUuk�փ�A��(��56���n[F8�<�uM�Gg�0��SD�8<�x�A�Iw �k)�H�8Yr��������/F�`FN����{ߗي\�0K�ۧ�3��O���Wr����o������%Ӯn������7�������v������W��J���6rY2���ںAO�mn��+�����"n{�1�ޮ�򞞬�©?7躕k�GaSÔ����gX��s/4�Eu����up]x����u�ֵ�t��,�Pȃ͑sϢ���esq��đ��[�U"K[20��"JA���D��#�y�p�,\?[����^�þ�*�J²$!$'o��I�z��֝_qsk['Z������V���a��G( \3Di�R�ڟ���zL�|ı�	}Cj���x��/�w�`S�I�怟��j֚� ۯ�QA�c���������q�k�uG�I�nX��^���!��{��d��{xQ	��C��E�l L��,��'@�f�'�\�^-����rB�������B���HX���A������<x��W��^�R���lEIX��P�?d�z*��e�tÉ��6v�����0a$�Y�o@#lb㹏xE��˒;��_�kh	�0�d�C��qAꈄ<Y�IJ��|���iǲ��*\K��v�[�q,�V��J�+��/�w��'�`�� w$�"��C�g~�M�����M�̦h�x�v�.ܪ@����5�,�3(/�(�|��#��Č�f��A��A <پ�e`��d�*��!����t��j"�J8����[�']�X��ێ%c�hs�G�n�M?���.l�#h8^Ej�i&�<�u�@ea�6�����]�i�"���J1%�0=��n�X�O@�������"���=���|z=�ox����+���vTST�h;` \�0!��1m�}�cmW7���S�xpk-��Op�{P[B��"�LYB0�A!5w���WȔ�Of�c�=����M��9�<��Wσ�T TY3�`���<��J�u��\\ �Ux)0�f�I���������_���rAG?������8�[ZR�l��݁�Z�_�� �9��S9��׊�KV�da8�%�	ҏ���DJ�NŹ�|�����M78�������"~��~}جα0���b��a=_���\eq��b��0��,L�0��O���Ǐ�����]�UDH#�o�a>�M��,��X̭�'A�{��E&G�Ir������9m|0�Ӕ<��������s�<d+Kވ~PZ��(��r����@<R(Ts4��I2v��n�%���B��=`��I���H�}zo!�p�#J�S�ޢ�7m"� �˃�5k�."$L�[=��p�#x&���1�	��	0H����O �$���my�WoPE���-���"JJwwJ*!) ]"�]�����~����~�'{�^k=��u���/jf�8J��N�q\�bO�'P_�!݈�����C1A�"v!P�,5��J(��=ǆ c��L 0I��y=����mh��S���x�Z�I"�'��\�z�U<��Rb���}����6t佫���IԩA��p�h�id�Ȩ�Bm�
����_ѣ!�~	m��B_4v�t��]Qz�bNذR��	('�l�xy55���?�O��2��ya�~�-`FHq�}�T�p�H��:&�E�� IY��Im�p�$�Eϧ�����#����*`�/#��LM�-���Ҹ\{�E�@ђP��=>�j��M��D���o��L��H����bIUN�8�:����ޡM^`�釛��@e��&�����WWR���Z�7�lP52�&2��,�_?cE�LZIw@A�@3���.��-��q��^]B%Q�ƙ3��H����~C�ꌆ�m�����6 �d60T��������_h�\7����ψ��K��j+�e��xk�����B2���n%3R+���:��:��R���1�����%��6�~�����6��+�����F���������\�C95#t�:G<��S���f\OaBe��I,�=k1�FJ�&?�Uv�S4�>�c�Ӣ��#$X
�d���0���썭��y!���4���3Lq��΅��
|�A��b��.����j�t���c�3��h��0mw`8�((�2iD%��)����t?1�G,�8
����:4�T%1p,�M��Tmu��)��˒��H������M�D3Ks����@W���ϻ8���ՔF|���H h��L�,������";@d�V�$�BXsj���YY(����,q�� �����})vr�gHaL*E|,���|�$��v��8L��
��lZ����p�B�R��<�����V�#�1,�L�`��0?�R��� �~�K����h������ժk��>봹[ֳI���}N)�R<!�ɳ�j���Üs(���i�V�7p��W����� �)��r���m�VM���c���Cuй��ot&�@ب����
�4���ĸ�x�&\,Q�t��.�*��� ��s7�@F)�g�#H�\x7�f��G��i}��ei4i��H�Y3F��X���e��7��'�UAP�w=�A?)��r+��/9L�ٴ=~��Ýҏ�%�^���xE���J�Π�-�����r��o�'� ��q'^}�ީ��b\�O�����LVZ�%�7$�&U٠s��q�p(�F����j݋� F�%���ߛ��b�"���<?AE,��B�0���� ��mc�IP8rU&ZVaL�����^o��9B�K����\qӱfL.fXF�UdR����S.f�{�<�$��$�Ɠ-v�T����*��q� 	��r9*�d} C$���kUeec��a��uҕ�^%qw�h�-������B5DM:�Wt'��}ŕ��a��ox�{��&ic�/��������(ȟ��X(h�&K����V����k�Y���X��x�6B�O=�o��B�H��и��Ջ�zc�ǆ�5:R1�ԛϬ���~�TT�s��B���/�o�Z���ź��5[|z6
s�bP,�d#0d��rA<�;��a���>r�}	���Aښ����犙�z� ۙ�-����`b]vn�!xc+�J0����k4�wA�GN��(�}�<x��̮�û�+u�.�X��ꕒ\���#TL+?��o#�%ʼ2��<iT��e�jp��Xl���+hX�����֖1'�W[�A�OI�fAHѻY�}��oOP] ���JX��w�7~��|�.���#l��*8���a��^�����'���J��<**ɷFV�Ӻ��x@V�p�o���{�9�j�l�	]���C�v�C�ްwǳ����i�f]���c���>Zo:�!NE�`�ot�@I#�N���]Z���4��K�{��ߙ�\(�͚� 3s1h���t9�t����ƕ��:M����T�"DN�&��j��n!��"��Y3�u�Ǽ4%�W����q �Hs �����8�Rb�/��nV��u��DtJ!���HW�B���<7��W��s ��ڣ���	]XW@���(q��i׵	\T`6vs�9<l���[i�����8�t����&]Q�S�b�+b�٨"��2���@�����}_j
Hc�||�p	2&]�^F�n��t�R���E+'s�8����轱w�s��Vo��7?������yjZ�S��A¢���m������T�*���1������'�C�X-�RΎ��|͹�tq-H�w�T ~��aʘ��<�n8�B8�� �'K��4 ������M��qY�}v�����_\Ұ�ҏߍt�Έ�de�g\O`�"�A��AVU���K���CF����VӞ���1���]��	�������=x#O�fY!B{��r�á꯵A����Ω�DI�a�z��� dnȔ^�|x9~�&��畘�1�b����It�l��c�Ϯ4�]��|�W檩� ��R������:�iu��A�O@O�ŝm�ϩB����9U>Gh9���b����-Aȶ֢��Pe�9[kQ}0S6��u��y�w[	��� f@�/��/�b�'�FV�u�G�(�h<]��}��)���?k��\�/���~ ��?�����v�7�n]�42�t���.O���w�4���3+��ԬUh�D7:0h}Cd�R3��Ar�Tcp�bvW����ć\�O�7>8K��}���"5>�Og�e@C5GD�P��趨�97s�(9�B7)%
	���T��0�F5��Nv|�`L%�s�I����?�mf�k��p)�И����~(����'r6������ �T7��-G��0��O6��e���`�O$�J'��Ɛ��х�K�(QS'�ͱ�*�m��WVg��,�Sr��w�<���TOK;�	:���*-:�?�}�G�ǋ�H���գ�-���&�������v�2����	jW�����&K�|��KI���IV)��d�<�$��>-�c�[���Ɲ�䱐���aMe��ɡe���؉Ӡ��D�_*��Ci�n��q#/$�dv�"�)#�8�W�6��їA��})�S:||8z$ldżYi�'u27�;��Ԣ�6��$�;�ԓ|0�B��a~\����l`�� ���YJ�lt�a�b���,:�r�qiǵG|���H�/a'M[�)��L8Ĩ�ze�{��B'�B�1{��lM���j��S��}�����_E�Wז� ��OK���@W/��z��'б�?hS�E��H��X������rA���9��3�Q��񯵞���zB/R@�E_�]`<��%�ʡ�����+'�WP�^KL\`���NC�s����ӟi�v��:,�-�g=�4n�Uk������������1,��덾	�Ũn+��q�Ql�ʌ��rP�Z��?�ݙ"4�r�e�w�.���xSn)y!f����ݻ}.��=����r��/i��H��c�n��)"$�1Hxn��������f���A����rZwbp��yw� c���1����Ǩ��M����nPE��K����{��s)(*���x�ɐ~����F�
9/���v����Y7WpFgA�̉C$��^��-���
Mh��CC�q��}@ F磗��a�L�[���^O�#ie2�r�DƜWd���QO�͝6j������3GoX�� &WKf��T'=ن�;�z4����E���n�}B@�1�絿�b(�7�qrі��ի�Js��5$I���q��a�ㅚ����?+qx���	eD����n�e,�B��܃d"�|T�#+	�]kgX���zQ<��&~ԍWϞJ&TQ��W�"Az%�s�É���CPp�:O�_sd�v`����U)$�wG����b��0�w~__+�%�W�*O-�=|
61�GF�|I?�k�QkFI&�Y;�����^3�/ݓ������U��U*͹�Y�K]�B���zN��/)*�{D���9.i���0D�C��8�w��h?{Q�*���7��Af�@���	 6��*3�H@_((��-B.&�/w8���K���r��w��t��~m�.�Xo=� ��%�ه^|� �Y�����c�՟�ؔ��|��HK��N�M�+-�=�Ӄw�����B���a�(�:\�/L(I�-B������D�W��N8Ҷ��]�䇜��I�B2{�K�G�����-�7	X��w61ĩ=9%��'���{�<���*�W+(��@�����
��0	�Sѯ'�+s��L��j���*{��O�g&��,)����(�-N�ޭ�)�l1}0E��gƒ��r)2�8�œ��K���>u6��q�Fҿ�5��?u���N�O��i����;� �3I����d�m��N����,BV)� �X&E�y��_ ?^�'M��=}��⭌y �}���*��x��-�&b��µcg���7�t%���g��96�2��?�'˷ �h�Z���E�U�%���>tH�G1j��2j�	��e�&7���f�4�XoN�Tt�z�h�GΣWeD}WɃ!)��:��JJ3ã!}�י����頼YIM�O}d�3 �S���s��[�\\��5���=�'��k��g1���Ϳ��u�q�3q1m��Vvغu0إø��F�h_e��I��"���1K�\Z���$ZG����S��TN$�]�C�םTj5�����J�Q�W@*%[�E�6�Z������[�\m�k>ʮ��dD*l�{�z>te!�A ������Xy49#�ة ��IL�!�����U����q��x��[w�Q�(��?�]�8�
�= #�y��3쫝ď�m��#��Mg�ؐê�d�3�/�f�ƺ�^�JNi=�H���%�� $�:�)H�����oձ��K\& J��p��CN��"�bM�&�
�T��d�g�{�3#R[�8�y���5�ݖ'�a���|�|D���2
�����{�453J��{8E:$t� mؑ��:4.��[tl��c �}0�e�8�y!��j��¥S������T��}���qi�'Bi�3�����,�z-Oæ�|Ԇ�N��,W����I���Y\�q�4�Je�XZAC +��KTqͱz[P��z�&�� ��:�;
b�d�&�D�'�D.3ǖ�Vhpp�?���cW��Ξ�+�ϵ��U��.���6dWX�z�m+�B��ڔn^^F��J�gY�~hy���1��M�٪�GN�w��o�X�a�W�Ǘ$v ����C��fpeP��b(�J�k�O���S�u�pTM���t�ͩ�F
�'%*��"qﵡ`�=W~G�ʓ��q��;z�ū�G�L����뗩�-��4>2;�h��`��������0�\���4nm�om�dL��H�&XH|��R�A�Ъ��RXlm~��"���7����DG��R���F��Xu�>$��'��� [���M�w{u!�\E��<�]ӑ��Bh�xe$mu�Le�.Q�z���J�a(�FD�����7�褂<C�N.��[�y��pZ�
K~�$꣟1p����oMm���O��Yz�UN�Y�۳�O��}��&7(rϥ?Qym�ᙛ�wO��̃@� �:r��`uZ6B^"VS���{�2����E���#�;ۗ�_�{v�$�jrm�����f��&���D�� �H�UMe�Eu�Y{(�OD��D¨گ2g�1���R=d�Rjj��;����m����!��1]͛Q��}��p"f� *�M�#q*\g49"݅~������Y"��Bh��^[�"��=�B
n��������yf�{$�a���X����Qe6�q�վ���������e<�:!& bJa[��x�*��a<|�4Q�L> ?��F���\���,S&���l�,/�^H	N��ϟN�]_}Ti�v���&�)���1��ㆉa��K\_�NJ�ĭ�S��~"I���|y�o���E�,piR?3��5��V�]3��w��%�3KJ����,0���$3������;T�$�*��w��j�@�=�h���g�)��-��bT5��OI�k�$�5��M�>�c7`T3��Xg��IP	������x����n6 �6�IM'XR��xԙ�^�I��JJm��l&���[���0��ؖ��p�����L~��vb�eQ��'�$��a�����4�b�D\Z��Wm~}8׹`�rq]Y����B`�4O�n߸��~��]¨ºȹ�)��c�>!f��:����5g7��7}ye��s��� �0����s�f�ҳ�ΐP��͛�v!@4\�<6�]Њ}O렫:���Q�r�u*Jfɸ0��mݟt�Z�a��#��KČ�%�;TYI�l�)�B"���Y��������kW�?�^g�ysT��	���M������n:#�溡n ��L��^1� �k������e���0_��w6����I�a�k8�JK�ei��U`����Tr������������m�q��ߏy��f�Rß$Ʊ�����������"� x��1���E|��V�)k�������� ��0�>W��;�ڼ�,k�\�wR�_���ԯ�XITmx ���Րde���*µ3Ocwd�7�߸a�~.��a����G��VK;���v���C����xo��9���Ŝ�,��MAZle�+���D��X��S)/R�83F�$~-�P�m�\��b˒�ڵ�hK뙥�ӧ<:�����8d`T�($�@@m ˾I�ȭ>��rl_��~�:|�g�f��jlT��_)R����N��u:��Ah�Z��e?U�����*����V�$��[�M4�
��RYV�;�Qe3̞~�r�?���?��f�CU���u�U����aH�¡�
?#N��r�8e��,%맿s�_C�n�,���_&��b���H��3%�%J�_mN� �7����f�N�ƒ_���,�?oǨ�|،�$��[��U�4��	Օ)z����KDDVFǧ��F�m`C��E����u3]( Jr([�V�s5�������7c<���r['��o5M_h��2�%.������Ƨ�MlN�����I��Ͱ)���
��.+�k^�8��s�nk����b\�L�o�}��� F����������������[?*�^�vV�I�y�'�+���D�	W�����-�V|��gF6a��M�}卆˓k��5�՝ؓ���'xD��u�'x���cհ�������t|l&_t�h~��G�'1���AJd$�t��q���.*�G���f�w����^x�1B|o��x�J�g��
���>�ή9w��>�����y�������(�\�;�{���F���5��O;�Q��iI�<��/��-��*�����}�|Ƴ���S9�r��Rǽ!r�飢�b`�Gp�Еl�C�L���#�o�z�fä�Q7��e��fbֺh��	x�Ǻ����]�@
0����>7iuD����Ր.�3uzoi��ϡh�Ф������V٭�B��B��T�����'ʤ��J�l�A��OUM#��P �-L�Y�z���p����r��ۥ�ئk����=B+����4^G��u�V��k���slh@y��,�
	K&�5�#U���L�	����ՋǞ��e�fέ�^yPt@�C�fm;��RwP���5\�E���	�ޯP+ˣ�jg�f!�:a�Gw�PBnƨ�~Mp]&&�a�d�F�"�l�[Q�`	:�F�ė��R�k��^�|�:��s>ٱq��1��շe��WK`��BIm`'Mv�Uװ��D�����	T���Y8
ٞ.�>��}g���WYV9R�.��P"76��Z�4%��	֣��a�DT��R]!����RG��i�����2s�KC���������9��|b�%A�7����xw���3\2��$u 2�G�o�_��
�	ĭ������S�W����t�q��I
j2��î��)�.����f�?���h�+i�|�Ϸ�y�&�yýE��keJ�\��o��e��t.zx���b^n'*S�S���p�c<�}o��̗W_?_����'�Kѣ=�� ٓ�x�r+����.)踩BM��%����5m~`O�g$�!~��	�ZP5j�I4�L��Wg#�Οu:8y�����e�����MB�i"-(>O����\7�z0�ÜM������􂀞1q��aL y��i��t�B�C�t�_8_z��ve�a#�d��w�v<~�t���'A�L��]z��.�V����܌0�`��NtcƎR:m�ǋ�B�e��o�<F��B�|x�zz�'��uM�"��������H�q����so8��y��]_G�;m���� 7]��#�n cؕ$�)�L�~�L(>Ul3�ǳ��g�/3��e�8������|�0���ޮ!��*�悇�.�b���C�r�P�a���IR( ��N(��IR��
�l�UAn±1^쁏1P�Ig"
���Ѐ�;�0�;�Y�)��EV3�Fb�䅍��f�- ��\J�˷hL��uW�tA}�y�iJ��5?�z$���؍�"���8{
����z�!��	�2`�CC��&S���?T03��~�e��Q��ڌ>�3��fr��&ǫ�l�yhρwɶna�\Q;H
�U��B�"�E�8=��b��s_H�[����~�L�L�y�1lh��������f h�gA?���1
I�A����|�����#��(�&iu�hP6�,ўWoh�{׆�עm]ߞ))�?:b0E�hV\ĝxv���~U�F�^��(�� x6�$Vf����%j�/�$h�6v���]���B�v�3"�W���o=t��8��/;Ң-��Ŭ��ڬ��ڸ�7ա+��� \[��F�z�a4�!&�dɲП�X_>��w�p8��z<_���%��f�� ���*�U������ݢ��K
K��
�N�o<����D�%C
KG�ͯ�K�?�<�=4i�n{";?|�d��Hh�Xp@�}>��^���n����ilp�U��V�5�j����{J�i������28�`����!��+���"�+���i��t#�v8���/�:�܀�l0����;kB��L>7@���#�Di�T�\UM�=S���,?�W�'��y���/���;A˸4�E��-{%PEUO��chp1���A�l'ĭ2G����7�a�>�����7�j�F��[C�d�S��n�.�������W�x�;O����	��OC�Ō	��x���ڟ@��	��&���m�=(-)��ʊ�f�^�骀m$� �g8�I|��kϱ+4�%��z�:2}
���u�}>7��D�Ȥa\&�Y�#5���	|�i���<u�|��Z�d���P�3�~urN��4�k�hBڪ�-v��W,��v3��L��	;��.��mcЙ= +Z�FU|�ߑ�Ժ�u�'��񉢟�qh�!a$�q�b�;P���FN����s��I��t�������`�%�A?��gG����.�oX��R��f��3���=GN�w��JX9a����h��sSYxl��fU��G��k��ĥ~�6a��-�*O�|���zq'���|�$�t��CS!C��g�n8�xa� ���l7�y�vjl'yY� _%NP�.-}Y��X�:O��A�u"S\���[��mh�&��GU��~�^�T���g��81��˒� �	G���]�^7M�
<^4��r*0lچ�,0�O7:����h�O>����4��ޭsQ�2�$f�\�8|� ?A/��^��ſ*3�XMA霫���J<$W���i�	�?��gOք�F��������lҠ^(S5f����l0�tXX���5}�̾L�3^�c}�"+,��AU�Wy��iK�5�-V�錆���a�r��B���i���؁W�td'& ��G5��'E�`B	�E<q0����,9T�CLY��O�jW�b��K��f�{\����>M�ni|Q�b
�ӱG^�J�W�s���fp����]i^q-���~oV^ܫ��K�(}��5�A0I�ڽ#���k_�Q��<��o.���tA7��Z-��hw��8ȃ)2qwG;�?9Ы�E]��g�>��˟��A��:�4㛘F��D�����		�|#�n��]Ҋ����oX��P�����H��{6�U��;Y����e0�sT�iV��0�ߥ4iI{�"������o-����tɸ�O���ܞ��k�#$ie��M��u^��A�!��ϱY��r�Vx��VRo{&�z�M�v�����әy,�!cZ�1v�C�.�G��S���}�����\`P���!'$�t��f�ȤaU�~��Ro��uAk"�j���7��A��_0�x�H���B�LĘ�A������po����V% w�s4��7��B	��"(GL���'�� c�3����~�*<�)
�H�.q@_��3҅�1z���8�$m������I;Z����w�����ڣ:~gg���S����cu�����@{Hq�n$ay5�4WF�~���(�(�5F�����l۠B ����`S�ƽ��}+��y��s��i(�ߥQ������p�[�@�:K3"�����Ս�/�V�U��X���4%$�'U�AH�뎸�?���*�����"�NϘo�z�����au��W��]GbI������@�+�Ey������d&Oʘ���A�$���Q�J6�Wߖ��(�;-�G��T�ڞMaq@~����[�n����p�b.���������g��K@�'j�8hLqq2�`j�T��FxhU���-��Z)���R$�p2M��<�QD���2'>wO]��^4�N4�Ov�v�9��n���n�5(��k6��:o{��aZ��C�U�8{r_<~.�3i�&��~��x��&]�",3���s:�SF˴��^C%P����k#��(k��A_)C�*6���e;r<�ϳ��s�:�'0�LS7�%.�.�XT
&9��	?�.\�>���6H�o؇���RHC���/��	�y��p�bF�,:5�A68>�$+�+eI���I�i|2��H7��X��		�9e2�_��PB�J$���m'� ���uk=�鷟Oy�RˏC4�_.rB�� �D��-���!Z}�d�Iy����}i��DŌ���œ�9��9J�T�tb`^"o%�)�"@�ǖ��⌵�tNM��a1���ʚq�*�����?�r>�DTF�ߚ��	��=O�[��5T1�C�뮻���B.Y��H�U�|-( M��f�/��ȏx��6H�����a��$�5i�ZS^S�� �	ix�.p��e��ƞZ8���a��F%��*]X�X��q-W�~X��`d� &��Ű�Xd��$M��C�jTQ��v�"���v�dGf1�,���**���d�#��?xH;��C�t���3w�9��#����Ԧ��gb�]y�����\�=�5� ��o	���eZa�"���K�o�Yh;��c�LG�PU��u�x׸38^D�:S|��P�|�����i�y��c�'����hb���v�B��2�)?�IW�$۔ı�u,�ǚ�z�GG12r��bΕH��Þ��Tț>�ur��b&��,\?����<yr�n��L~WR;a�b�)��#�t��Oq�b<�bHb��E��F:�0 g_��R�Eӽ5�������d���m��~4{�����Y֒/&�Y9� �\���Zh����Qe8o7]�31MF�1B�8h�C`�ʙA��!�'�9�����#
g�Z5@\%ʈT��%p�OM��f����9� y�"���F����o��̕_�A6MJ�"4�zz����No.����jҝp��H��1���'���Bݎ���\#0㒬���3�f�r�c�������ݧ�'-ZEm1x�8��Ì�����7��J��3X$Ӕ�jŰSE.����%�;�+3_��+��e��Y|�L4����7qh��kr �~�s�ȵ�|�5��&LM@�����&�ԥ'T�!oL���E��#M:�E��]���\�u����&㊠7��[H
F���*�1�lV���ʴbQtc���%
798ҵ�̈́M��R��E�m�K�� S�ӯu.*� E.Y�ݙ_H�GS`e�\p���O��*�E=�?PM6�MG�n���](�@)���0�ܖ��|J[j�.�;`�;|;�(�#VJ��� ��g`�p	{�0c��ʥ+~Hn��{R} VՑ
��g��HI��[(�4��ٚ\)�Ż~��?�Z�!�v4ց⫿�y΁�-c�v?._���Q�i��-x<���yV��}�4�L�ȿ���d��7%w|��䃯���$��4�����<u�<y�ŻYk��M{-��l�"�
Cww@P��Z�GHH�l�m��:oI*�Ed�Ou�8P��!W���q�������ߢ=1���`��]C0���x��������^Q���MG\�>�&#�A֔q���1���{jV��b�6B��4`�nn�ut�<��'\�?�4>�`	S���4��/f�,vzc�����'\���� 뚙(���a1���L�T�����>�
�Sr�Z�
�˟�$�f`X �^s�8=k���JyiJ�r���(R-@���I��7��۲��bt��,ZB���g�*�{�X��Bw�{�G���r<�i��1��OS{��N�D�G��r�k���H� Q����r�F���Z��ϋ#��<�(�	Eۛ&K�/.�4�YV�����a&U'�t��F�eؗ;g*��#+/p��~�>�������%����~	X \{�F��C��X ����������ɛ$6%	���+��ټUx�=,����=�L�;~5)Q|C�,I����{w#�w�-���n��t�����K�9�7)!����^�$�|l�b�1�w��I�������'����v)n� 
~`97���fU���~v��[�@(�>bM������]���;���w����yj���$S�6A��v�):�R�@~M?�q���t����� ��V"��-��P��qǼAr��V &��	vQ(�����Tz�ӡ��G�x2��b��X$� G�e��L+Ѧ%٫����9���y�R�ь��>�A�(�aa�Q�]^Y��a�[�Q�_�\��F�0>(O���l�����0>�:ݮڞ��>`���O�JJC����O�	�x��j�/���ښ���&��D|U8A b��7��%�������KlYvoa/������(��Ԁו�p��ED�x���.�і)9wb�A�� ��տ>�P.Y��T�T����͏����؟4���_h��DX	rP��X?�:�,��X��m�
���%��������Dt� ����eS%$T*�~Lϸ����� ��%� C}���$|��A ������,N�N:_r�Oۏ��I�:��[w�~��_n�8/�J���ȷćP�%;l�Rih�'0���	Ü�)~<����Ї�Z�u��[�>߸���x�``(�n�����#�:f�7+���4�E�t|>ߡ�"l4p�����P������nk=Չ���&��%��`ʒ7�����=�;��{�3"�x��h����:F�����W|���$TT�(
��0Y�'�����ʯ��P��x@)���A&�����9���|���D`؄�rֽ�]6�8��lv���MX��cx�����r_A�糰ߌ�"���aq�13�;#�����o+�Z:ӭcڭ�}L�m���mUlq��w�A�n�K�i��C�iM
�?+����?t)u@����X�ot��&������J��-؀�����C��G�nt�����7z���7�"� ��T�|%3��^|8}�=�4u2c���9N��cB���b�,-߿�����J��3Ƭ���oY�<&vV�V��l�Ϸ�-!��D��|!�3)=�r�;͇}�"!6mq���mB�!��R}����U�N�a��P|Q�Ɋtd�g����`ZKR���r�h�F�$:Hn�VF΂Dppt^)�V�H���x���|-]�$����]p~��2#�&�Lz1m1�g3����L��f��t^�;��?:�"?��D����9��j���y�W��I�v+��1ďlx�������`~+��|�;���FA8ڪ����+�dFo��9>��ɶ���5��|ۧ��'>�%c��ǰA_���@�|6�Am-H�*ߐ;WTJ�(��D	�֬X&�PXQ�!�������c��U)��᭣#)��`:K�&��`^
�P��ŕ��|x�m�	h�G>�2��������3G-�|�\������K�O@�}P�U�^�Zm"�@�;>G�ok������U��蝧	{�y|����^�-��*��9M./�
uh���O�S^|dYE�Pgw0Tu#Mu+���a�U@�/$�������|�kjҽ^�,Ӻ�{�~��q �8oP�����x��E^�+
ʻ� |�/����U��0�s=��UT�Ђ����).�/�/pM���r���V�O���nҡ��I�]��С��g�gޛ��җk�]�3wr���b��O��B�'�\R�$'���ߘ�ԋ�$�\B����-t.Vz�ս��0i��^b7w�µ�li��jPHN�ޗ�sĄ���F��|h5�e�-%�a��p ���<V)�(,�in���	G�dKdyDrX<O�c�j?�D�}�������dVuiξ�n���8��ji�A��S��f����Z=���h)��� Y���[P�E������Om7�W^ե��u�>z�.B�|��oJ��[�W�I4_��[Ci��^6�JC��X��pqq��52�@�/<$�Zw~[���&s��H�R�����}�A;�������iܥ��L��[ �������
�D �_U���FB<~\���r�K��:��-��
ȗΆ�����nx��Q_-��T����RJF�����=������|��Wiz��q���$G�?A���*F{1��\��O�ӧ0��@5D��q�-�}U6�R�gC���Fr	�
�7�C�Zt=�c��G�R��p���P� �����w��ڭ�S� ��~4%�g��!���"ĪXP�[�}���hZ��ĻZ|�����pH��<�!{\��&���NYfygQg�Ay�9VI^����S�� �C�.�Ǖ� ��[�pF���;F �-bC���u2����]?�}Uf`U��j�.T@�kP����@���oҎd����OeHO�@���>��ra��-�u�����"T��k�	iߓ�2����\:�.����rU؋g?��+$����W<�+�4�d���sf
L�����2(�aQ���&nG#��ަ�E�Xͧ$p�P/����c��A����R�����ݯ���������lB	�,��\�NW��_=�?i���Z�c�`�O���f�gUD �X�W�2m'!x#�����P+y*�L�����0�~��HF��7r?!����֚�C�ö��5�4��Υw4vuX׽w��P?рX��u�&� P���0������?]���y��pF�6��i�֐do4�N���I������a�S/4��A���p��U4��,�Q����]S}�!hg�s.���>�
ɋ�Uȅ�ϲ�(�!�\>��e���\"N��'�*���s(�sy� H Xz=���Oِ��!�@����>	���Y���<AX$2v��.B�!��	���S���@�1�%��>oA�C�V����b�9���.�HS�a�Q�������"	�9�U��X�7*���A�h��Rc�U4��TB/6y�8�?��F���� ���1<2��D�" ���C�����ϟz�-D999����:e�J�o�����pZ�C�����Ӌ�8::�??z�0��c�w546�H��Z��
�KH�mm����jhhdee0002��=)�q?~�rnpS-�r{:��jyҹ���Ï���ef֪P���b�j�2��g�;���9��.�'^�|~qѵ���~j$)-����b��Ι����	��4v�@�t��FFN��8֮��o*�|fjj䌡�Ҵ]�Ɉ��t�q��b���L��'U���e<NtX�`ۥƎ���g��Z/��{�N4�z�F����HH]�E�l��2��SH$$$\�?'��?���e


L�e��oƿc5���XZj��QSS�?�e+�ozj�TPՀ�(�r0-��m�,��f�e�Ԫ����=�N��!�m�|���2O<>�v����7CSV<V�iƄ�D���$&]��@��/,�����������Q�A�O�}}}�O_�}�m�"\j�F�p}d��ˆ����I���%���LИ�Э�c�̯�6�G*N���e/�d�ZkC0� 4M��s�=H���B�QPR�|�����!��=��wN˯ IysuՃk(SkΊ'iaaQ���be�\�yڒ��}���ň��X�\7��P��n}S��9��2����r�¡S8.�v��s���SI⼐�`w:����I�ߚ�������s����4�t�������<�ys�+2=?l�0�d1}�@+��p��x��j:�x�����lYI6�
�I��Y��##��BvY���سcf�=�9"�8���z~���v;�u^�q]������n�����,+���~h�����}�w�4]����G0kM�9�O�D$�Xd�[M��jk%�V�5�1�599J���Hy/���C]�nT|����"�[��l���.�Q����=<44�eX�hu<U�f=U=�]l��P�f��W�Ҋ���'����x�Ls���߹�I(9C։�3z��"}�r�9i� {^GW�G�Fo�"��g��go]��P��[/E<v^��ƛ�y���4�2K��Y'�h3[�u��R��<�����M4rҮE�޽���U��m����7���-���{�����@VN��`{bp�Qjq@��\԰5A�h����=*�Ђ������(�R#�,55�N�2�Xii��t�$��-�W�V�,���.&�c�Q���<\��f�Ђ9�K�_�Р�TVm�{�n�S�Gee�PԆ�S�������ڦiFg	�2�����]��R`N�ii�jjj��߼y���s�Z��������E�st<i�zz�j`���TUU)��D����I�7-��K�����K���|%o��,�B[W��ĸ����0H�t����e� ��tVY���� �	E��$A|[ݨN�����̽2q��@(9�	2�:�jc�����h��T���(eΖ�W���^1����kll,;����}�S5�J���7��ztO����TE�&�l&����l՛�=��~��
C�Y##�� Τ�y�����CPP���;2*����m�<���� :j��m2������ tc�S^�lDN��b- �@+�Q���$�J���/�b@/�.�ʣ���a.1))��#�o����9
�
B�m���]�n������N�L����.�D���Y&��o��;+،��IE@8v.���K>�L{�^��G0�����7�}�Y ��L����|��]�����#O=�n���6#��w#���~�f���0�5�ɘ��H 5��9��`�����z���޿��o�2��e��u�~B2��+|�܋��.�gqD�*B|ngo+��<Z���Ջ�뻎����/6��є��6X9[ĶwdD�`w���t=u����xu��d1i9˿�+�š��iA"�VZ��l�>��ލ����VKK���h$���s>�A�[����ܗk0���_jf�<�~���3��ҩx���ǟ����h��Ј�"~�C�ti��o?+,{������{�K�*�=�R�H��:��{��Gˣ�w��f���P����:p�Ժ���S^������(}vqq�]��8�k)�6�K�A1���i�O4:�A��S����V=%��~2�t����U�c=��a�o��-g��*6|%][��Z=��;��]4��]-��J�v�U�Q�v�ZoR�}MQ�s߳�?��A��;�]p��j����P��h��rF���& �m�-�,L�d�d%&������DQ�۹�Q\�G
yL�'��@$F����]���-�뉙��i�̵�.��*���Sn*�n�y�{�w�/ql� r&����&�)��2�GA���O�DE�f*6�)A��1��r��8��������6?���k�<�)�P表�h)oC��D$�7Z�����ٔ�RI�o�R�-F���bÚ�jaz{��f[ޫ��kVr�ns6��>��Sc�V-��yѩ����'�^}�_�^E�?��o�������9��� �l,J����8�40���nPf�����%݌~���ƪ�}؂�)�h����l�踆��t���t5�]LNO��g����ͳ����^of��E��]}�����뷦�,�w��Z��盛p���6,�҆�1��dx)�7�־�rZ���t�R8B���Q|R����������>mb�Q�roqH�l�yX�=Y�+ZYg�����W�]���$�׿��vب{��M�D��c�a�蠟���	d08�ggg��K�LC����n����
ѡ�(fc�gye��+(X]kEQ+F�>;�������F��!�e���>���������_������NuD��6��9��e�#�ݩ�?K��X�i+1�t�Ň��*��ѪP��+���o��`�
�X�;6B�]�|v�L#{����P���[<�x�b8��%.M��6�aҧ�1���C��:L�W�c��	��B�]�L�շoߞ�?.6����Ȕ@��s�`zr��?>�����$�ZKJJ����p0�)`�֓��=���(������W_0B��$�5�����#��� H��3���e0���}�}�:^����9~����eMsP�#P��M(j�޼}���ic ��dc��9�~d<�T�|%MUM-�<�����	��8?�꾝���������l��B?�xy��,�]�-8Z�,K6k�h?a��o>��#�����?MAR
$�=�>�Z���]���+EgP����Xg>��MJ������3��Y�Ǐ>s@C�wz�QL������)\��a|�0��w��M��:�_yDULZ3bhr�����Z'eeR��zR w����"��8������vc��@���^�,wF�'�������VT��#>�*��Ɔ��J� ��?A�GM~����"�J**�;��LN�!l�

ĉ�	M:�n�C�a�gx�h� P�Mw&��J���7���W���ţ������{��"���1�Ŕ�F��y��W>��>5[Cyq$��H.��5���z_��z1|� �(�Sj��؎7�iVQR
��)�ӭ����'�0�?�y��{ڮ&�̭�xGZ������33��v��W�Q�)W�q;+w#��F��K��t��$!�:�'O.g��7:w�	���}a�_Q��>������72r/7��4����,4��� ���C��.����U���1d����)D �h?/[ͱ ��ɷ�����f�g7��oE��ݴ������~EHHu00?84t�USd�n+`�}����'G��&B>���.����L���M�(\�����[�	���-�������Xa�x{Ր:^��hQ�Y�EO{O��� ��8-�<�~�5���o��cz�F7�֒���t���D�� Y�覆I,����y�����O`��# п�$%%���k�h����"�7���̪��ɹ0a����ES9����۷oAh<��0r���#��`�c�03jM��K
a�O�����LU�q�|�[]__Q'�n��;���	䢐�@'`�2�cǰ�Ǻl�PQ�!��������L��:<�N��!��~q���#�:|�I�?ߌ΄�@�U!O[i=�%O8Ռ�mzILd��	��#��A���ü�<))����X����N%��Yw���y�z*�i�ګkto��2T�ߵX��	��!�s`�r�(AbA�Td����*_��dE�`�	����������6�����K�~�w��M �H�v0���A9>iO,����)�TE(J9�X���沲�ۗŢ"����98�			Q.-5i�_o2z�:*#P���	���0b��>�
=O}X<S9�&}�֭�iB[��8�`������׵�2��7�`���=���>H��;��3�c�GևX`}̄飦E��9�����3��C�l9�C�SSS9�K�S* ��t_���FK8%7'�(������j����F��R��T��_F����'������pG/�q����$����2`c؎��k��fBөٱ77[��},��w���韶ї��S"��T���+�9v�m<�!w�l�!��)��*�;K�t������1iT%����l/T�l���^%�`�.�.�3i�o�ld�����`��;�a�t�$$V��K�||��8
M������a�����1����<f'"
X�I�f�Ws.�A4��k2���Dy`���ɽ���(zW\,�
��MK@#3 �]�U@M��=y���:~JJ���ѿ��]AG^�L�&�l�x)��&#�P4H�`�{:4R�W4�K�~Y�'&��
����-��E�B-�Kdd|bV�]".�����q̈́�7o�t�j@�8��ƖX\j7Q�;��or D�8O�+��##O��hM�y�iX�h�յ5�~My��{3�����.9���Q	�- 6�4��[y/�dy�!��\��8P�@�Š����}�#��Z��=�5��8�o׷���7N[����8
g^�~-  Mև.[%桷Q����o�B��h&	y�%�Kއ[�/�Ύw��t�x�W��,ux�0W.� `(v.�8\Y�YK�����L�L��MP����>qa�|�M���[�XUEV�p̀����$��C�9���^�� ��	�c&���'kI&Q�1b�ь���K�aـ�=f��ɮ]�Vd��!`P���Wc�F(�w'����C������������ ��4S�z�98$D�*�.���0���G����V)GQK���H�b�z�EqW�]k��W���Wj�	��#��҉��J��Jk�2���u�]������s4 d�:&%k�fqi������ϒ�F����a�ٺ[`/�g��޿j�k����(r��w@F�?=,���K$T����hI%~888X�J��5euբ3q��%%��l��G��o&�p	�Ö~��(j�U�n����X>�����,6���n5G�Ha�c��wj�S�6�1d#�;�A���׏mm�Ë^}���#���t�F�B�S�q�3k�k�pԭ�ULn@bJ��P�5nͲ���	 ����G�nl0!���=z��A~�ڵ>9P��z����{dv8O[l܌P��&M��u��x�`����<�0	xy^�|�-��ޟ?�uQϑ��o���U:�yB�D�U��^���c�]�;�������oz��������?t�?�,��;�g��)��U�_�]���f��%&͂`���[������9���I�*Y��u�^/L���%�:;ǆ%z����)�����/�t9?F�4����'����fvG3�cE�@��f�26v|�*�w|����6=����� �'�W*ڂ<l%c3��uAZeK �ꑜ\�vc�Ңrr��@�9dT���Qs���[댈�zڎ�SE�NIc�����	u?����Uz3�V�Xe�7��������,�u�E����KVcΏ�MVX�=�/p��bV�s��/Y��ZWb�?�6�("""j=0��� �G�(���_iQϽ�s˾��ư��*h��B��O��M?�g�	���:�骷p��y9��FW܊��}�骫bV}���&� T�O�~��t-鞀 ���3m�B��_Ш>���u�G6/��}n�x����kY�@�}q�AQ�1߬b�B4�G��U��g	�ɫW65rEZ����`ev��v&������H�B(���Էn��x5��f�n���4ѓ�1����vNٳ�D{�ژ�	r�cxs�&Չ���Xve�۴��ь��p�8X㇘��d�9������˶N _G�7���	�|��EN��/t�E��w��B����BW��D�9�_�N۱�a���ɓ��6y��h�4�uA^�j��?��]���gprr��U���A�PC��>���@��ʎ���Vl @�4�+)--�*�Y밠=55�4�NPP>��mIZ`�O��rCI�뒱:٢̍���$$<-��Y(hX���P��@ZD���r�P3�����;;hI�~R���oh�>�ׄ��Ԙ��.)K������H!aO��4�[��ɝ��.�i��Ȏ0J�.���_g�ޭ��.��W9��}W$k Oֻ#��n���q@Zڟ*!�#_7uth�� ��!�d� � ^3�5ϫfƵr��%A�bzh/<-g�G_�������ŵ5���̀��qAq�@@f���N ���9�}�z�3�����c���H�������Hu�3<_n�J�3���`��"U�y����v��?�g�z����!o� \���[R53���'�&���0���dy�X����]{�$��FzGW4�e�	�f���U��֡fi��HrQ%߃!�el�S2��q����m��W��LJN��y�jզ*�c��ol.p; ��m= J�C�fUKBDz#��p�ױ�����#Q���	�v<�f!qV��Om�|�@�g�-������x�&���wI������/��/�!���=CͶ���1��Y<>�`�ZT ���)�iH����P7�~�{����5�)����8��������p��������m���{��.M@#�"A�RRQQL��Ysrr2:ٝ(`�u� ��B�T�E�_�'�����%�Tq��� �P��lE'�?���f�+�M8M�}�jJy�p���wwz,yEo�+�ŋ�^!5쏑���:3�.Z�PSSS�6ke+/ c�b�;����	���w����D��c��H
F�����Z������� ��<0�5�L7�|e�߿6(Ohx�p�� f6���:o�w��W�����_��r�\''� h�KK�e���(M�Bn��T�| \��d��:��q�
.m:+�����!##3|YY9]��ff} <	
���x*��X�_�&�}3bK�#�pgie��uA���%������$��AP��f���h��m��Y�����z���O@��9n&�����cjzX�7���|� �0�zBQ�S��x�l��p�gWF��+k� �)::;����W�~��͢�Ñzw;�~����]8≇G�P��`�޹���X�˸n! ��d���#e����ȝ�QD�i�ѓgJ�;�@ ��K��Kn����P�x��L��Q���P�jy��]Ґ?}�����	$,e���2����i,�4������<�G5���/�l��C'�4�o��ʰC��)W��?h&�s�F(A����)ތ�g0���B(��h�;�����C��K���~/PѢ��g66�;�_A�x� r�x��I�7G�:�\4�;���dDoQ�ů?E������㑬,w&����
5=����$��	�rrr�1�.+�S~���Q�ªϟ?�OE�`�]����*����S�vJOpߤA=�����"�R��;�q{�I��m3�(��
z�vr�����	%,�tyg]h����CE=�m�z��)��qK����߲5�(.�-1n��F��4^�`P�ħWb
���ӧ�}��O��{�gy��U��J��m�Oᓔ����j�~��~'mmb�����^Q��Hͩ��":��MS�١� ��˲Rm]��3��((-*"wqq�+=�=��@����||o�O5U��pjN祶��	��+Ï���_�����Z|����Q�/�����P��#�ti��u�����fUs��>�� `Y��z���@u=��[�'�tٴ��w�Y��������&��yVkZ_[�Ρz����jI��Mw%ZV�J8)�r��;���ЇN�~mZ��s{2�?�.@Ҙ��'�^���>z��"��?~]]�_مu	,S�*Ć2E�:���44\����ꐗ���
�Ͽj�%���E��_���Tmʃ#�zBa��J9��0,Q��o���d�ѹY[����LZ�,����y��b��,��w�wd��˻Y�Ӯ�~N������4`�$`է���!�o�AW�����)0��I�/驩�\��r3?p�F\T��/�zlG�P>�[̌$�.$D�)wjQ<�7e����$������pk����p�R�����U�������ӋM8,�n�����0�L��c�Ǐ
��_���ܷtј���������0�;�ʤ���xܱ9��+�����B�&��I��yP����5����(�r)U�!����Y@i5x��_�/��ђ�
Q����;4"�i��ک7���uy�c����D�o���kA%�5a�x��;UBM�'"<� ��%�̔�T���< !ttu�?�3��p����YT���|�ɚ���|��D�dI��!�����E�C`�|1��.6`sE������FkO�!�W�^����S�#&{��gymb�����5��Y�������wŽ�͕��6�B.�WӤܺ1�F�����G�k�I.��{���9�ʄW�ù���t��Pt�u��x2��!����Z>UU����u�m�g��;é����!.����5�mx���L2�F���fi�(���|7MҥmI|�W\�x�w���;��{,b�5��V·PQ67��	��G;S6c�	���[��>�y�t�X�l���,��+� fzv��� �����������kff��6  K� �wU�a�jY�_�PMX0��g��p>�j��n7|��	EP�C�ߩ�0�%,ﲄ�����
���6�7Q ~�gk�@����5��bFj�W=��"�)�
B�u��r��j�A{8v��Smdl,X�[]����]w�@QGF��x��L�[Nr�v�R6Y�ѢjP)�g:"n�O7������u��@�	�Y�'������8�&F����
����&�%tS&䚏�xycg	�����E�n�|�[��E���C�m[�r���������U�MUG�s�����{��N˙�����&*f�� S�v�������\ 7�q9���p�Z���$�y���P��Z���pq��Eyf�V�N𵍛�먭�nG=q�-�t��vh��W먎�1����O�'�E�563 
�^JB�k�̍iϑL����kq��r,+�1�^7��T���21,3%"'B�)Y���oX�xciz0 ���&�/H����5SV�J�%��Ϳ�d������w��x?�"�wV�� �V8�H9��1�ͣ�g_�� Sx	&������]҅u�W�)@.Ξ�5�j���==��G(L�O�=nu�@'�y#999�%N��m�gl��������
iWO��#���� ������l�d��:[�B�K�0A�<"7����*���N#aw(��|'�cM�$>>%�CLB]�����E!S��{���;v��l��߿�DAQ`�5h,+��S/՞`��XW����kk'��O�88���~~f�l ��=��8՜A��Tv�/��'L�=V�n@�5I��r<SS��Z�౷��v���%�����o�������ʹ,�9<D�D3I$�Ny|�:񭜹z�*���eF�g�T�]>y'�n �����4:�M6K�۲�����s��<[ɞL�@XE�H˧�=^-�3��S3��6oa	�Z	��bbb,����ru�M�_������:�K�pr��nlh� ����n�c	���^Z*�9��Vlp��K���R��ŗl��g�9Rn� h���MgzS׏ �w��4x�ǀzv=����v�1n1�rg�yV~:^���y���M���M�mc��l�p>k��"����N�˙�R0���J9O0Ɍ���e�ӌ�2D�CwLQT
��CD�4��bl��
<-m���}�fҼ�hk�ov�5�-�n;�����Ņ�$<^����NM�p��~�HP�f�sՒ,fԞ>�:�u�1�:�ۣ���~���6J	�Ch�#�E��cV/���C��i��gc����6o`(�j$�sM}�%!��l�/hş�xA�%��F����i$�[�r���wGtV�&�d�����[���;&��_�b1خ�+��o��5@����5\<<�G�蛑3��t���q��)yyվ�p�]m�_�e��r�ӥ��q�ᅔU �hD�;t��`����V���	 1��X,J�<a�������O�=9�}zU�M~p'`,�N��)�ε�%�|��f��A3�� :d7t��)G�-�+#6	����>���cb�Q�}�����H�� ��T�(��*�& ;�iii��.�nGW���s뗙~��Á��g�r��,��1��X�e����6�(s��̄/_�D��t]��of��_hj�:L�n�Qh�R#��G�-X�� 5�bxѫr@�E��A����8����zujf�0;N�H�E������w���Pb�e���C�$���5냙�OLL���#���ױ<
E/�Q5��D.�ب�5�i�S��k8�.�d<w�5��@7�� :D{���m@������W�OUwRg�B�09I�⢩��u�����{�jB`�13y�L{ �S������T��_���:�a*�pt<�L��Ԇ�||j��q��`G��xQ��H��w|�]�S�A��:����yyUw��j ���7����~�Z�Y�����e򘆖V��"IQU���徝8Y�6��[��:�y�o��=Bb�W:��;��y_P�����ifg�]�G���vI��E9���AJ������>��$/'��\~�����x<k���(��!�Ϊ�#ׅ�@��H��6��i�w���ؾ������gk��.����Eޙo4,2n4�&t������jia�uLCU5�s�=ҾQ�#�pb-�=�@�{��v�r f���z�vJ��U�GDPK8�
o������@g}�EE�߇l��/^|~��^\�	,����*5����N4�>��vi3��*��G�_��X���� �h��Q�p��l^a``X���E�v�"������g���E'�Of��G��N%�h�����,�le:�o���-,,d}�3�#���FFF兠۱D!��f�5�3@��Vs��eI?��H����v��; %&͎5����S�48{�&˙���ًH(��ݚ�����|���L`�4��κ���s��@��\��s���K���=�w�Ė'���~[?<�a�zsH�Ð'�iLJ?t�)��������s���T%T��n����(��ϙ3 P-Ȫ0k}�bY�{�'~B������E0��?����W�#�+��B��So�v�=�	R�x|jj�����- G7���OO���^Ɏ��}��<��D&����}�2����$�-3�u��_�!w�Q,��ݹ���B�L�be!غ�{�L��G���E@&��&{��A��w?<�'s������z�^S[ww�wy���T�a��1[�����p����2/�;�Q��2��÷�}��C��-�G���O
��85�������졩d���)8�
(�@�_��:��W���x�۩�`!7���r��?o8���X�����&�_��Q��&Ss*��6�4,��_V��R�@�h?�$]ǚK:��ب^�V4�݉?^(=�6cf�%�|YU�/>5�o�ى�
�q\�	B|�:���m�f��m:ojGhC��Ԍ���tː�3���Y��w=
"��	���1&_~���{�i*�f�"9��b�.��CE�b���`����$�,�y��Gu���^�::8x���������&ج=�l��lsɗ"nj՟��]F�I__���F�Wn=����ɫ�C-�\�iK ��T%����͛� �8L�`�X�(O޾�U#6.�ߎ%%sP-?��������*N��݆���� ���ܟ�����s		!�փ��Kzܫ���1P̐�1i�e�����lkV+����w�D%�|�0111��E���ح�R����#T����`0��e�ſ~�89=ep���P66������v�w�($?�_��B,�k���;�ߔ�r�?�>VU�͜U�D���::�ƴ�s�v���ttU.��6���U���8?5��Rm�����J��J��\����=�=��*t.�V	��;;u~�k|��U��������I�g�y����˟g���~�:���y�}{����l_�s���6�Ѥ��T��h6�-�| ��or�qn��`0h����͡�4�ʜ��E���l2?���&����Ɉ`�O�|&�q�^[�G�]A��W�>�VB�F6��4&v���`��϶|�b
U��O�|U�K.,?�>^j�{)��}t��w��e��bs8�%��:ۻ���g>���w��o%��	?�k������=>l��Z�>n����r�#&���{g��~��_;�]Q��ͻ��P�f�4KQFaF�FLZ���%�Ʀײ�/ZL�]頏�2���ʍ���po�ǂ�XB��t-�@K��:�
�ji1W:� W�)c�������o���/*����)-5y���~�7�-�ԇ><S9��:�59��uye{���{za
o"��u����s�R�9���3W�n1����i݂��ek_�|�p�
�O%����9������>�(&���f8���p٢AʖQ9�y�Q�2&;f4���N	}�w��P^W�es)�5��l]U*S�q�ƺ�~:�S�������>2���z�ǜGk#��fk8����1����X���q��I�xߛ�{�Z����c��[��o�t྽
XS��4}S^�m�T���pLy��fR('a� ��x A��pB��1�h�ZpO�ږ^��T��o�)a�1��uwǬ����E�.Cx�0B��#5���I%/8JV��t\.%$;�ҷ�e��}@@߅�>�P*Q0��� PK   DU�Xǐ]zd� K� /   images/700e9707-92a2-49ec-8e41-72cbd6a28b0b.png<zUT\���n����6xp'�C� �� 	'��4hpw�����ǽ���sN��N����]�j�WW���I�	  p�e4  �������u��Bp��$���< h
2��^&'�h�����*kE�g3"��n2'�5�k���}��z��k��Qr*��zQ�E���P�AU.%}�����	�;ޓ�k�EA�������5��Y����� w�+H�UhQ`�����	�dC��_'$�Hn���o�)B�х���Զ!b�`�[�������߰5��:�r�v��khL �t/�����v��K_-)��i7�8yol&�ө�������;�FF;����d�^#��D�a��|�����i�2���O,i�B�K)����SJ���	�d�`�-ǺU.��I���_�a+^��G�+�X�Ǹ��K/R>2��W8G��R�%�.��*ou�G��/�H�9u��{<i��'�G���'�*KR���k��n3V �6\�;l̊�n��K��x9���r���9�/�J�h�~В,y�t��J����L��H"ˊ��r�k\�}ff�ƟgVH�a�
�q�,T�l_V]z��)���<�#=�B�6f�z!�]&�5��.;ޤ��V�������r�{�n���������)Y�km��~��$�� �gz�����̸YN�#�f��x��~z:ٞs�t4hӨC|rS�ǅ�9?�UFr��?M�?����|�>\�5En�$GF]��O�=�_-;���>|֧=�!�����X�38x߹�s����SǮlћ���ۂW"K��� �r)��pﺐ�9��_��vw���ֶ�NW�Η��G�ZVe��?����Qۅu��|E�켙Qz����̮�+N{�%��U�ݪ͚D��L���Z"k��Ǆ�J��%�k���< �z1�*���Jy��DͶ|Z��1��3��
�ٴ�d7��[�7�s��y�j�sL�kH�\�o���H8��t:�5<�+#��6?̮>`�H��&)ο�P111�WwN��ڧ���*$0&}h���:%��d��d��۱�5���a쳨*����'�A!�+��G3�)�t��]E�0G�4|�@�����]�=�'n
3ާ�����0c�oi�-3g_����Y��8;q�t������Bt1pVc9#⣙�tӷu��p&��������(w6>�T��i�
��i�|4��@k�lHش?m�J���敒9DX�\N�(�
<B��T0�+k�.e���3��	��!���*���l������Fυ���w�o�Yz�]O���)3��P� �������Y�E��a�k���VUq��in(��L1q=�5��s��,'{1��L~ ��d���<m�t��n#���y5��ξȸe�N<�B�x�h���0M�}��]�C����4�|�ʯ�;~�\���<"1F��0���(����cCgK���;cqC�d�����5IZ�ln���_�Q�����Wnr����Y"�ٞ=�%���������g�)~-�����O���%ȈA�����cRdR�}t � bn�����8U����d��>��i�����IN�_?!�}Â)�ӃfN�j��z��{	�E/�vj�-��gBrh���F��FX��AꜾ��h���G��I[�l�Dds��if+�Ṳ�q��>�l^kE/ݧe��>��߀e����·\\�������<�!���GPeG']4��k����F����?TE-ݐ<8'k+s�0��Ш�����x]j��U`C����]�D������/��M�'��⚊�y��26\U���~@
ش�+K�S��CZ[w��`n\���p�A�u��h�x��fcƷ��_�c��N��!/���*~G���Le�Aċ��
2����!"�0m�Oq�ّ��o�v��'���=�r�1Fحt�i��BC���يO��]sB����n��@����1��VМ��K(�}������	�}�(��V���%t�p��UI'�^�P�7-��K}�:>bk������Z�S�W��T��sW9}���}#�>�~�����Q�bР���bBt�rF��Z%~2�c�����������B�!
ؙ��μ��pu�S��Ɏ�PF��Yۅ=�5�[�e�J�$����sC�(�"�tc��2'v����%�A$d�9�z�����w�TmE��꽍#�)LP-��>#��W�.vw6=D���
	~ �l��"�n=w����p���Q��Q,��j��LK�7�vU�6ϔKX����{�����3fݥ�VH�����W�+�s�ȵ_G���fz�+L7�e�8�n.�Ґ5�2���#Λ�N&-�Y�P8�CC�g��|-:_,��{���4�zb�Ð���Qң��P���I xP��� �@��pR�=�� �Pm�3��|��l�Qd��5чV���A0�}�v�{wS�� ��jX �)�s�e��"E�"�����kF��/Oi{ �n�*$�<氿>�O��4Hg_!1�fc�U�8�c��ke�R�9)y�(�6N��T0�tUi�ܜv��]�e5씪�ٓ�f��%��,�b���Ǝ��/CJ����zd�(���!=����*$�G�kq߄;����s�r� �QZ�V��]��zE-s9��8���ɛi��侮��չ'~�A�s3�TU�����#�(�G)�-�K�=�m	�S��S5u����U�ܮ��T�}[n{���H-�Yc���~�ը��{�����=����\�����3B-����RNB��_i�J���8v;*k��g�ܶ[����AU;F�$]���2��.dA`�� s�w��8h���~��x�~?Z@�뚸��\.�pD��O�����h`���@��X�~J��K����|O�_�᩻&i�1d��>[�7�:�1�6]�bW�RC�E|6"4|���l�tn�#]��u��J���o������a5��/����o�{���-i�{nu]W�; �z<	���_��(�֫���F��nM��d0��۵�@ ����ˁ�2�v�t�Oܦ|k)>��+4� ��=��o�/�%��~���[�92��/]/{N�ק��}���ވ�&���jwP
��dm(�AN���z8����%�Q�Aܕ�����@�/�U�s��D���gK��N�����WL�G��un���!���O�U��f6�2�*�?`�
ui����^�q�*_���ٷ� n1M�	O�����Y�|^[��~�R���_1�~��~��|�;��bP���"�g��訬��b3,{tt��� �O^)1aw���rнvZ�q� Jʗ�)�5�+0�n��y�4$�5���Ga`�Y���H
e�5F����~<��Z����s[�a?����̴�P�^{���>�r4�]��f�+�l��1�tߖ��o�W�{q�����0�Eد�?�$E����.��;w5�R,8'T	�?qepF��zf�!�UX.�i]Ͷ��S�/N��{i�����Ǎ�����sEc�7Za	����B�	O͐�Ւ����=<J����fE���s*�U���2�
�'�N0���ߝ���m���A��՝~���~���ߢ~M��ņi��j��LŊ�k��x���f��{�s|s��Κ&�K�-z�$/�g~���T�5~*�+�gr	����>a�܉b�*��M�J=�Ӊ~��^�7)z�f_��$�����5������o)�Fp�MQ��N�B���u/<��ڬ:z���='��?���J&�:��8����U%���� Oc1c]�O�z�h�/��LŶ7�h�\!�~�7)�II����"�����S����y�J�M�`���]�m�MN{�xh���Z�s��ƚ�u�������/�D�r��s�2�`S�s�7c�>�	ճ�'�}S����Ӥ$�����J���WLV�����5��t�����K���x����q�kd8U��4�?��?�O��¦�T��_�L�:�,W�^��l��H`T�3��P7d���3�����(��"����N(^��S�Q���+�K��������⼋�Ѓ%��	�y�9����݉���~�}oܴ�&k�;\$rw�J�`S�����A�ۯ'�u��n�|^ú巏�㧳n�k`�'��S6fV�x�M��� �����v0�ړ���*"�9��
ٸ_��`n���9x~ �e������\o��:���7�%&^���k�?�,܉V/�B~���Ia�3�q�=N ��t���=������-�dU�w�$c%���>~���O����c�)�#�O��4���w^�H�R��I�Jq7�@a�E*o��u"�E�F�L����̬m���M~���;��J���S0HiJ�2���lB���b�����OW�Lfz�g��T�m��ԏ��	������-����;��Ґ�(H�I`�.[�%���(�<Pr��8F�"01��>�/T�PCS�:�b���(x��[?��I�������_��5O�)����� �=�m7��H�y���c!#�Xm�p�P7<`��EPD�����Cm�?!���[1�.��^���l����p�6� px:v�ⱡ'8T�,���r	��X?b�@��@��&:�̛�L�*�׹��4�J�e$=�{�
:~|g����|�!������:N��$a+�9������*Z����j[
Kg�����}Eze�j�lM������B�Ϝ*�I�@=��6�/�N���D�W5m�}0�� {a���W�q=?eHP`9�!�����VQ�?����*rJ9�q`O,��L�H�����������K�ݱER�a��@r�ȴy��P^H��`P_��u�������I�U��bD@?.��^�Mv�wN��n�p���[��a,� ���B]X5���?�qzP����I���m�wcK�lE��5���OYh�,e:+���靏b�HA�^eo���ybW5X�9��YBޑ��T�Sb��{ni��z�p_
R�o�4pc����i�Z,����`v�d
ėbv�W�!�4�wj�N�*���y���3�A���[�/��&���fX�d�oC4�
���+2Z�B��$R���
 YSu��P��G��L�m�*�+���mVp�]V�ix��%`�/�]E�-"�w��M��< V�7�ȣYL��k0�P�g#��ڌ������`~o4�c�0q#Y.�4z�������e��� $4����㪙��f��zǕF�S6E�)�+T"?�Sq�P�ߚ�(��l�j�����{��w_W  ����K�ru���-!fjm��18��="K����ڿ���Q������k�uFDgD���?j�KmTk$J��	α �X�����$5�1,7��~�����d��]k�����)p�\�n��.������F�{�jƎF�d̴���mX�dvg8�����3WHC__!�ԫ�[��[�	B+>E�2��@��3h��5���'��f�}J���zF���6>/M�9�ϝ��^M��b����[�j9��9-��*����Uʥ�+M�J�m�l�U���&��7�䢺����P�b&�.��_�1�N�y�>\�z�9.[	���ǫ�K�<�����Im��:�m��?�+#'?Q���ǟ� �J��OXgv�>���{9��=/q%l��C�f�:n9�*)&]��'�j�LNz!Xkd�&me�<Ԉa�J���O'��O@��4h�wL���ZYխ��xQ�C3�.#QT��R���ٚ\3	\Ԥ���ے(�����_�h�
��}c���U��]�_���Zj~�jr2eec+��d�B�:B���I��^�$I�#� �N��0�fe�q��gOT�U6���� �f��]ۑ���}\���b����:o��ɗ���fb���\�茆�ژ!��Y�x�������P��?8����nch�i"���շP�Άh�'eP{��̻����{8i�wa^�b�qw�vt gls~n�����@�7�JƸգH�_!�����t3�V��Ȏ��T���|������� $ ��r!�8����Y�X��;�7�2W"*���+]�Ի���2������o�P%����C���ҍO���6v��V�)�	����X�$��w�<�l�/�}��h2ǟ����ӛ}�K���	��Ҷ���]�(Wgf������Ѓ�	�zmmu�%T(����F�sY1n�O�+hb$�$Yon�w\2��Y0��r�9������=m��������h$���Ğ+}���ǭk�z�Y��Y�+Ĺ&5P:���H`�%r�|��%�sݛ�t�gw�i㊗��]S�t�B�A�g^M@�'��@T^$�_�l� �x8=�"=M���w�%Z�2�Y/��O۩�'u�:V�2�U8֊���c�v��C[Y���:����0�����Xшo_�������Q��<���Lhܦ$ad�{&���w��E�<��*�!H�u�|�^��M%AH��7gk�8��%{�� �o�̸�)�����	��O�	���	����)���@�����A��A��kD��>�t�m �D��8�A*�m&e�J���<��c��U�I�p'<��]�+�Y.ܤp+����MB��~���=�cN�3�������m\�lkB����W]�ǩ�P`ӼC�gЈVֽ�&���b��p��.�<ߟa�/ۣ�6a� q�L�o�A�L�^t��y~��e���������?B���:��?#;
_NS4{��/)N׫��Sl�f�'M�2�X����<!���ݻ�{�F�W���n�'6՟�����6�̤N��t1h����e�j���^�d�"r`xC=By��K��L|?s�����卟�h�xPuR��r�}��nc�0;Y�m�	!8�A����&���O�ߜ�)x��!2�:������=���7{P-h����bШ�h@41+��	`���}4WF�I��k�!WhS�L���}�9��"v�[��m���Q�6IU�m�gY\CT���ǥ�ĬG�)B�Gs-�D%���єj7������/>a��/�:��uA��
��Y�3`%��Rc_�x�3{��d�Щ�r��p�i�XV,�L�ڨ.�[�n�r0TS���$�'�x�����]�	O��w�\v!�FFDx�^�͂l���|X&N��3���P��^|��؅��:ϑ�\ ������ �Yq���-����q��C�J�z�@�7�+&mk<�e0��~��t!�b.�OY����R�[̘z��p�&}RUm/��ҿh���ߟ��/I��_p3$��#��Z��&'p���ɴz��o�s"�X2�)q��z"O�)�.GP��X)m_+����'G�u*Tŝ�kHҭ��.�mȶ�nX
�gg�P|���,�%:i�.�"����i ���3��qS�W����4�R� �v���esCd�~��w�.��u"�=s��bv�NC�  �s�0e��h��˙g�h�� ���8x*���Ծ	���R׊�5��᭦�{1g�jֿ����_�{�Ǥ'lRc�z�#0-���Q�4�41~��-���)��.��������jFZ}RJuq�L�*`G����Ҫ�Վ���r�J���9�ի�h�������m)b�/u��.�<��6��2�BM��-������s�O���U���~��͙/�dyd-����[�Kq�mXM{Z�/�] 52�"�T��-f�\����J�k�V�k���U ��C88/u�H�Ġ�@��y��n�/��(�Hq�"���ȗY��ea1B�4lOeu�g�kJ����s��͡�8��"�5D�{�����+05�L>M@��Dy�e�l�I
�ȶzw�����A�����a��{o	�=@U'���Sd�^�����ytz_�_����u>̷Iw��mћ��܅
�l9O�sF�����|5�:���	{V豝�A9Z]Pg�{��~�C�Ƴ*������1����3!��(>��S<WcQ+q��c�վ.Cy�qP4.�x��ǈeh^qU��w��Ƀ�a�rN�d\�%�3�D��]��	� �4��fv��E�c��6�^1E��v�	��_�
�@���r��l~��h��{�Ag RP�~'�r��p���1*�W-�/
�(<Ȅ�ʐ~�Bu�켓� ��hx'S��A��6;F�q6�E��>տ�fUZd?z� ���H�E�9,�GE��S��$]/�Wd]z�{��¹��Ju�1�|�9>���U#��E�����?��R!v��%�
ٜ
�hE�"n�漱����5T�-�ٖم�ݮ,)J�ܨ:n��$�A����h������vK��z�GS��+&�J)������z�H�T-�Dج�4��3�LN9�u��`�y�
�>^P<�I&7��/��%:��F#���oɒ#N氎��d�۹Zs>o&�4�#�'A���)�f�*���#<�Ͷ�m�w����?d[���8��ƻ�U�ET��L6�J�D�:go����&��[����(�� �D�E����7�y�P��;�Ks��kn�m�*��r[Q�Q�"dH� ՙ��t�_2*(�:��z�n���B�Qi�N-�;B}�ژ� l0ZVnD)���
ǐ�2����[�;[�E�E�,D�Õr��,�%ܸUx%��&�H��:�e굉������'#�X<�7B2�����R����K�Xoo��&,�T�1(s�<�hM������+W!R�g.:�O���";#o�~ˎ���a<\�{�iP��ś��<3;�:�=��nzg8l�aC8%Z�*�ŠÂ���o�����4�&�·��X�*�㢶B����츉�˧��lo�a:�3 ����T�;�)w��C������R������y���Wg����.�n�&<�u�^���rr���zȕk�8�|S���/�� <�w�L�Y�;ӛZL�)D���k�V�����\������]�I��ӹ0a�t(��\�j!̾��\�x�?�G�i1d�T+(K�<I�,�i��w}���k&G&���P%�D�Z	��5˘�����g4c�<�۔c�;0)S&�K�;�����<���Q��ϻ��ZTt�]j��J���l�}|��\��UC�y�Z[�Kժ!�E�Xhucw4%\2#"Al|��ƀժ�.{���q�L�/E.TC�oI�Z�x�b:UQ�1�!�)�5����DšR�*��_�z��$[�)���M��1n������cbP��4��
h�����V��"ǜ�?}Ǜ���߷ߨb���Ԇ)#���j/�����ٹ.��>�����t����Ƌ���M��V$k։�$[8�#�7YYX�z��q�n��L��Ɵ��.�?��>B���s�8l\ϧX���ZBb�$�]�8T�nLm��'|~?�ʝ�K�����-��������u[�X�6�Y����[��K�m�$)��Ȧ[�'��c��cɬ8f�7A�W^�|��p����?"�WՈ[I�$�2�w3s��a.Xl�u���CPl鍍�[���͂Lf�����Px�Z�������;�4<q(m�o����+��%�w����:T��=�9J�4�[v���@M���Z�<+��#	�Y�\gzj���;��%W�7���v���Z�����gaG
&��o������uo��\�*�Ci�Sd�齅�X�K�x]~�k[Ä�������pa8��'���;����J]`�}pF�$k�aӿ�]�b&j��ZHJ����[�Nj[��{u{����m�s���N�Y��&ݙ��qw���x�2�Ѭ)��W���g1`KzI�-nzX���_N���-�#�?7j`��r�/[�D���\>�u��L�Z�13�o�B�9.���h�4�$i2Y���"�����,C�؉Υ�-"� ����u��p���ꢁ���g@�������۱�`�=I;���&j"����NmJ��am٢�2WP�&gr��#�2�D<j H�(W���B=]��?���Nf����/N;t�"���t�}�tOF`��S�+jRԸ���d��G�����i�H$= %Z�}u{c	M�0];RJzD�<S���u�v�Q~)gʎ`B$��Hf!��+Ֆ^���̠���_=��8ABL���Bq��zb���R�W�rImK��� �WpK �=��c��I$��3��	�Q��_���z5ʥ�4辉@�:,J��'&bY�A`�xr�s��sm�hD�&�+9�O����tk����q����Wr��`~��� X`������֛KS��������������)��ő�x/eV�C+,v� ���*S��yW��<~ �4� ?�$�i�C���V��w��`�����Ub�`������Y�%��}	H6��P����B,"�G6��xW�C����'x�H�T�����e��W�<7T�GN�����'[�caE~Ks�3�JGN��t9���3M�_Ռ�-�y�;o�S�������zC�c"k�%���6� �b�e��x\#�� �q�|��9�s�]��eM�fV�E�/��ą?&s��:U%0Q	e���F'�ڇ��U';�C:+��wބyMy����*Y��|ǫU{L�e�,�9e&�n��«4h�&�4Rݴ��&�K�N.�%�Z2����\،�z4G����lk/V�E��e�s;�
U�����du�`g�sҾ�$�9	\�������beJ�P;ߣ�aml�P�y[�#��������_�a� ��ƶ�s���� ���n�
��	���nҠYD�OY�aM����y���u���>��f<ݽ	N��Y�&�����eq���{���9O����(���&~M�� �Ѓ!��?����*��!Ѷ#��!Q����V�C,H6�7���0]���ϭh�h�c��9���{N����?�����h� �z:57Bb�Dy�D_%�8HB���Ys���ęS[JsY���@A��O�^&�9�+�k���e��(�n߹De!*���-�a��58��:�C�~��p�fiF�1�1�1Cn�������DJ�m!лTWN'�,����8�>���A�
1����c��񥧧��f2����e��I��������"���=��!�� H���=c����rj��,����|6m۰�8!\˱��Zo$�;G9����mmy�cm�^�QgHTxIƕ���N�8	����˭�Uܐ=�N�>le>�|�i�̀�ާtt�x�7�u�<�o�es���"C5>��h�c1"Vo�l|M*��q��wk`Q /-���$�y�w1�@�����Y+��]w/+�� ,��s�׺5)�}5~T�a��i�o��hH����?�b6;���OL��5�|C�i7X�<��Ϩ��<���+?7�kao�`D�)@Խ�ː��l�?׿��G��_֎�A�PAD��Hj�#-��-�xi��3 �'�H�H�Y�-�"b6�y9@��=��zW�A[O����P{f�)���*¯h����3�B٦_)�4/�E2m	?�M2�h�#d♍�L3�����G�7㏕2P~.�3N	E����������ܝ�B�y����yO�TA��z�/&���BP�d���u�;`v_7]|B�I�]8��Xn�2h�87�{݀�%�]#��;�����ʈ�0bA�� ����#i�a���D}?Gћ*ɻ>q4_j��^q!��?n8x;WR�@!o��(��B�Z��hh���_�|��§r�/Y�(\���i|���S#M��5��O#m�@} 
ܠ���E5�������'x��\���'�y��̅y�Ɠ�ѧ��d�>��*���&�Q��tI�_1���3�`;������B(�:Y�P��`�<[�NŘ#Ή(��op��Ѥ�y��M�M%�j�w�Xۘ7֬`����R,���/Uk��0z��?���wD�0�V�~i>�"���/W�S[�?V�DHBzs!��5�(v����\������fDh�PG �������xۙ�����
�WR�+�j ����x�Tt��p/�$���������ĉ��;	j���j �⎸���ƊweI����	��k�X�13�\��ݓ}�
�_w_�����=���HO��m�v-�S�-�U���8I�N�����Ln�
ɭ�s\d�ɸi��`;`�Y[�Gji��ґ5�*��o�!�C��)�������p��a�z�Jز^%ʔ� �� �.��;�X�I�Q`�G
�y*�xf�3B��C��@���%"�<>ܜ���7��MƮ��b]���o�m₌O�<�A�@�g�Z.�u1z�����D�΍�u�S�fo2-���I^�R��t��0��M����8����H��h�ff�8��<�M���"v��Tؠ���f�����z�՘C��Dٟ�xɡ�oe�����paRD��W��1m�����* �k��<�.� �wo��.+03�W���[���bUQ�g��,����T����џ��l�-�+P�	�x�Ar1ЀBc��1���ˏ�wJ�� p�oN9+:@���8��RKbBN7�N+ӿ�crrO��[�=.�w��d(/fj�lV��&X�;�ϱ��ຉ±��@�;�D3Y�bCY�L�)��@Pa��6*�S��[d=#�["���R74�����&�֦$I��1S�d��[7�;t�]t�^��7B ����q��u�N0,KS�\�X�(�8��C�q14�*!�B�^Ϧ�������ę^I�~\,ߦ�Sǀ |,l���[��!��z��[ɲ��JS2��Ԩ���L�x�����6>	;�cYX�S,od�HK�0�i��ᓎ���o�m�Z/�ӻO-f�U�F�c�7m�����	����;YXj�̓(�$���H17���x�ӻG�.��Y_y�vv�	�tww���mrTRFq�+ι��nY�tj�?Ŗ���uY�{砑y�o��6�1��"��5�7#��1Yʴ�	��ϙL�x��+Q��&+��Z���Y�=�3�֖q�K]�*:I�����$!���t�Z(q�oXI�jdB]t�0 "ÛKΊQ߅��	jɐ�>�!Tz���}b�d)�`3�]��m�Łs\��=��=��e��m슧ў�  ��vM��*�Jҧ���'C�y\F��F�*?r9;�uM��I -v��R?Zy�">�IY�s�ʍR�=�-A�<�?ݓ���)�P��vX����{��1x̤j��Z�c&��O��{�j ��c>�4wp����Db�w]~��"�;j4�^��r7W���t:�0@����;y�o�/�xzX«��J�3b�v?�
��Q�^n���8��8  �y作���5H�TT��\U��XNym�3�����k~��ƏwC��J�H�Ny����|�l᪑)�=����'V������ ��^7cI�ǧ#[e��̜�O���!98p� ���欕�`eF��E�Y��z���b7�(�)���1Ż������ԥ�~4�� ��$21{P�[��_=��V_8�������%����#
����b�����3?��.�Ow@�^���H��t�޶��/L
dW���_��I�:��J�.pG�}��`�eQ~3>�/��A���:Y9��a��5q�Lpr��;&U�a�6*����.����a.C	��u�ջ"$3"0�2F Y(.R�^*��;��+�E�h�|��7϶��]-��\y5Iư,O��2F5���"oڶ����P�/����=Ah>�j%��9��
ճ�����T�����C1�31�w����L!�����
l�ɚ&��s��c����R��D�<RS��:�wc������W}�Z�ꊲ�ȁ��>���T���1_�~�w�Db��޹A�v!<TA�,^<E��BF�>ZX5�k�~Cd�Y$�
wÎs
f��&��@v���v��s�� �:�+�Β��,��yw�5�xr��G�a*+.�pZ:�B��/�?"��Ⱥ�F�ۋI�,���xs(�0_J�v��;W�3w�-Y��\����������Opr�Ao����5�čM+�ѯ׵�P�^�i|�puc��VϪ� gd���������-�9��ɗU��0|Co+�b�o�2Avn��ʱ�H�$p���5�w?Ұ�����+�
%3�B�q\i�>�8�@��ꒈ�q��G�N�sYA��5�(�"�Hy��l��Dc������9�b����>b&fT��Ȧ2�C �(��g�	�
%�$�襒��QU��Sد
���K[�a���p(2�gr1 (��z�=�9�Ш��&�H��D1�������-��(�".�ءF�� ˋ�و��S�W�P��������m��N����<u��Wu�x����H��S8D�܏�q�;f6�4�v��հ�uA��%�4%5H"���= y�1���������*����Eo\���uә����I�F4�"�#b�k���,��g�f6?�;U}�j{-�W�� /	�x�P�nĠ�
��n'�+���\J��OQ���q$"��$�S�J�8ƳD���C�. ~�o��$8F#��/r>󞆫�ſ�A��>E�~K�;���&����Q�ꛡ?hq_�~&s$�V��Y�|Q%u�i�B��hM0ۆ��"/Ɛ�O�'=��Եa�I����J�������e��%�ҀH���EM��,/S�?�D���O'�AO��g�h˔4�A�\����Y�b�:'͎����'Lc~�3^�D���G_�����$�v�OC��-�����?���@]"��J��<��A�����q�Ue)s	p�HbԽ��w>Wćf�/�u`�JA[w�o��u�����4�%�#�4�.�RJg�-\/��g�Q��{�|�gTN��[�)�
�MҫA�9	���c�W�zӎڽq'�E;HG01���-���+p{
6$����Wo�:��MF���fv��f�4»Őh!�s�g�A�p�IL���c-u�N�����)X'k�ȖYQ�N����7������7��B���R0z��	�:�8F�o���ԕ�)��keO��ӱ�MV�S>po�/M�J��mJ	(U�ӎi�V�A P�N_i{ �H!A����s�;ć_t<!��ƥJ�3��_.�$����E��:����s>�S��<��+��)�/Ma��{qX�1���e���ڧ��G���.S�>&j"��~[�´L��onYu�n˺SG�0����jG_����+��#����ی��N��t�9����X����k���g�ĳU�we,�ڥ��tM�ӾV�{;+ks`�h�K	?��[�U"u��#| z>6m�}��z�]������)��ltĉ�O��I+t\ac&_W���4��-U/cO�pܜ��U���J��ݸog#=��s�Bh-�(�TyuyS�@��{����BES�l0�9OBPqO�B?���5Kh�n�3��B��Ry���ѴX	�
/���w�VB��"��SY�e���t�8'�UG�I��W
ζ��H������#v%3*�k}n�coO�j�g�*ptTN��"n,�W4_��;bª80������[�D\�$�:��Q0����S w"i�x������]������X�-um �}Ko�P�b7�~�3QY6U���P�z��R����<�U� �)\/K��w�L[}1A��9JM����y����=3������_,�[�#�w�Lm��H�wEiV�8W^	;�2�ն�GN臚f��a�>��(چ	�������'���r��~��I?++����<K>j���O�B}iW&�ڶo)$�|�4�۩�;Š)dc�!�j}�vs����W�U2�=܋$ooL��4��+TΡ,݇eC���|Į�:k�5�I�?���Q��o�� ��ٯi�������g�u�&��՝���cL4���{ն��.n��Z�P�䉨�$�P��vzK�r�D�%��U�f�=�Ps�~0H�?�ԙY�����Ȝ>��#|nh3u)�'u\ד3lr̽��g�n�Z~k� �mrXWtߤg�0�xH�z�w;�7)�+ pIJ��: �e�ypG��޽OI׫�H�\(�'���Ua�S9L����] ��J�o@��
]'��ꊆ��Ǐ�b-D9��~�)
쯝!�D�XM�o�����`o� �b_K�_��=�������NQ/�ڰ��ķ�T*�WS�0�s� |@���Q��T�kTJ�$Tcq�?�����=����S9�Z]�[Ə�����?q�.�%����?�Dwǎ�裏&#�p�F�(_Ck֖R�����9ulv>?��Dh�J*�ї��VBy��>8k��2�N�|���5sf�|���>ӊ�U�.�� >f�u�LW^y9u�O3N��2�F| �"5�a�z��gì7H55u��2������?�T���/���������C�a��.����A��.a�ʕ�F�U����w�Ü�
t�Q���ߓ���./��t�J���~��ʶ�;s?�0d�զA���=���1*�#�1�
�����i(p����������ߗ�)e��c��~�q*-]Cy>����0��Ր�)�z�L�8�y�B���T�R��ǐ��<p5)�*���i��/����P߾}��4z��_��W<�x���P���V]�VZ�t%�0 w�o}M	D3��`fa��ul�[_���<�\�p�$����@�^�CѰJ#��B��Q��������~���|�̥р�}��%ũ���f�z��<��^�֮[Eu5���ϟO�7m���uDF-/�D�FO��/���n]����x�*����Abp|>8v�}�������$(���|p�Y����}��E�6��үi�UL[yL/��w�U�6��y�Q$lq�#p��}z�,Rn����䂿��Rԃ/�U�v��m�/嬟�d-� 6e%b��E�ԱS<�
��x+u�`�r��d�9_�IlH���?�<��xz	�q�i�����oyQ@>T��.@\ȁ	��W]u;s�>7��i�TX؅/YĻ$�#%+��d�jJZ^ڶ��:u)�+����� m޴�����iM��j��ch�"|��5k֌��%%	�*/���ϙ	����M�\{���*]J��EG~F�֮-�Ꚑ]l9@U�:*[W�Lⴶ���4�P�+;Ā���9�1 ��G ���'��'�� �����6��;Z��m��+)T���nZK�C����p�x�h��-4w�����A�!CQ�>�U������j���z���?����W��Fz�����30(���ѣa�E�xS80�z|A2<�o��CǮ�.�3y��(�08�4=L��,�mٲ�����8�^�o�2oPC���1�%�/�0��0 ��\D��y�ƏF�:���ҕ|m���(&-_��j됴.E��A���N��������իv�m]�w N��JQ����W��9�|n޴�^{�E:��)�>Y�a-{ư!(�e�__���	�-���#���C�zı���]���.��
P���JgMǃ���Ac�r�F�֮YF��WR,VE>R�&ȃt��o�<o���~D�5	��۱�0�#0aT4���j�.��K=�#����?�����G���V��+nG��䥗�kdz�s�"�t�T[g�דφU[Q��8�$�[n���)�{��٠[YY�.\��Q�F��(���о�m]t�>˖|I��7?[�N�hU�reo���D�)Z���o;ڴ1D	�K7�p+���y�>���|��t�L?�}l�#p�WΙ9�QW�Ϡ}�G�z�^}�?�����)�{��tđ�r����5�LD�A�QUU-���@���ʫh�I� h�>�(h�6<�r�<��s,y�a��T�38��sU,AL��+3n A^���i$��IR<
�~,~���h���޼�i{e�?����O�K��u�_�=�Ye.@q�Yԛ�C���#x�k��o��ϋ��a;�@:��Q�1��ø��&�
GԾ}7�2�H�D=���6�����2k�!ھ}���;��4v�g�}�����w� u�������|����u�d]s�5�[زq=�{�%<�7u+�H�W,���6;�;*�%h�7�(�C�_������^�3N��y�OӺ5k�8�����r��!�Z?�Pv.��%]L�J����?��:��R�n;U�l�bҜ���i�hݺ
*��Fյ�}ޅ����{���w����d�>x�W^y��}��!0����@rA��u����LI�C��6�	~�@�$D�'�Q�C�(C�> ���K��oSUu��� !=:\���7�J$��������i�?�۴v��'N؟ƌ:H��'b�1�<�����d�Cy��dz�9:���q��H��g猷�z+��C�5ft������4�#���nc��*�B���4�d"BK����D-�UUo�H���>�c	2� ���Bk�ld�m�Y���I��'�y��ѳ�=G���6� ��Fh�$ZG��O��舩G�9g�I5U���I2'�u�z�Ek(/_��HY^
��Q����P^�*9�l�!�4�����p}��]v�et�����T^^��@;�� " ��. �C܋#�2�[층C��WD
zUvB����:� =OЖ���ʸ�����S�~�bfgVt�_�>�Y�q��i��8��<�ݾ��:w�gy�5T1o@����H$T1x�l�k�Oe��y�*� �:�;�<*�ѝz�!��1���#/8}`�=��C.L��O<��:�(���5�T^V��!�����C��C�E/-Y���7�8�|ew�i���胏?�pK��>�x�6��7��ɼQ<�d�w��t�Yg�AÆP,RK�U[��r��8"Q+�d�^Г0�F��H�G�������/���x 9^��	��#!�����R��X���D����M�雯>���j
�}*7�O���─px|D^?8��L���c��/W�w�t_��8`��7�?%���[����U�D�Y!Ês�GdL�rN/x���ٷ� α��T��OU�CN}�ʉ9��g_PM5损~��0�í;|�P'��|0���do���v��`��F�j�����G��W�i�F�rĀM6�~��!�P��9�D����#�������z�x���4���l�>`�lauG�M�<�N;�T�ٳ;��VQ2���3G������CAC8�î۷��	�@�g�[(��u xб#�� T]�u��JE/|�����2�2В�g���i���H�8}-��y��L��iS����T����={��h���>�d�@8)�'ڎ�$H�I�'6��Y�(��2qm��R�Cg$�|�53i�hX�6�PR{�N���R�G���<<�˚�W�ʕ��r]�̰XK��
l�f<�D�Ka�+m�}%�0�2&^)�g��� ��&��NU��ţ!WOD� n��#*�ߏ$��j:��{��, &g�M ��eRׂB:��cXY�=��Gh^)hc�n������!�O;�:u*u�܁�-�џ��L��s���^�U�V����`�׏��Z�1���i᢯�w��[���1��T �G��:��?�A,���S�$vk����*C�eu��WL�,��փ����C��q��m�����x[��o� F�!���oLd�|����|�s޹��c�q�8 �A0 J&����^ �-^�m߾�>s��d\mg�yLQ���@ｿ��a$*A�i���z��co����D{x�n���[��7��&/��A[�L}�	���:�Sg� Ε8e�Ef�.y�)�+I�dao0�C�����p�ް�����"�8O���[{ђ�幄�D�ޭ �,��G�^Y�2�������	��l#3J�F����R; ���<d�a�MR^~'�<�p�/Š(�|\���\1̲8h�w��s�,��j�5���!+�|�|��ǻ�5d�`���0)�>E��	�1�H�_,`�eH�P�����4�7��G��)� �	w�ѣG�ĉӞ8�M�3�H�~�U�Ѕ�ϋ��%D"|=p}��G��(�+��������.��w���3�������z&h��iC�J%��1�DurMP?y�v�F�;�S��Kp��xRe�D\��bٚ�����Y`c����r_�/�#�s�^��8�3W|'Z����8�8Ydd!�׽+�,���@�%ͷ$��;��v�eW�FԂ'�+�"���) �c��[v���󥾄 ��&� iJ�E@[ȿԻ@_�x����kQ�I�O�w�}��_J>3E�D2�>#)�� %y����Qu�h;�б�<� ��GT��~��ڸ��~w�oc+�?��G��]��c��ǜ9s�D��_"��%0����!�"E�eG�>GL�E�@�{,ؒ.�	��
������vR"w�ഖ�6����$��a0 �m�F� gܸ���v���D͐ÿ�b��z+}�����/2^���g��#G�y�����Z��cၫ'4�>"�ҧioJQ�f;��B�(�f?�R���������>��:�*����ۧ��L�j�}t�Z�P�|�  �F.�s�'1r�}��/@+�X��~�i�jc�$x�#�
-����E��sJ2.NyN]C籱�H�~�|J�|�� ��� ���Y}7%�,��]zۤo�|��ޘ빂�|?�To��c���CGR
	�L"V� �RA��ku�\@E�=9
�5}�"N��r���!��&v����O�;�z ����pA�0�y睼c�Dh3�;�v��(�`d�1[�h>X� �ʐ���?\XTpe��i%�������a�hDe~T@Z�dᓉ*�������<0T&����@�2R�"�
�P���q�����s��>���O*߾��"���@����j�"ڼ���*D�f�Fzo�'�d�챐��Ճ���k���K�]c�	}&�4�
`�J&�l�dLu�_^�e�B�H�Ut@����:��6�_�r�����
l��,$2�B�0�E��.� Y�t�^��m���N�Rr�>)D$�+�Q��Y(	}.I���`G����+�0hp�	����G�+���@G�7pu+�G^�H!/��F�n�����;v�	����{��x�ͷ�G�|���#.�����v����(ʉ,��C��O�%d ���� �%��HLͿ�c�\�^�I&\&���ŕ�`�֪��)��,&%2�q����ė��q�G�|��CI�!�i��G�d��8�A2RaZ�v)�Z��k��^Z�v͝�1��*�����5�\ku�d��'ͽ+%� @���g�E ����`ӵ^L^	�G_bl�ѩI�����'=d_
wX�s�w𿠦p}�nF�`<ڀk�}E9�3
 $���e"�c�w�L�_��SG��<�h�����˞���~�/���P�}w����x�V1�Ȅ�X��=���~4��IdQs!Y[�s�X�9p�>���y�F�����@�����[hђ��������@�z!�3(]��t-� n������@d�q�$�t�v?��

��5k��m��9mz��U���f��(���D��\�.����f��Ź�q��`�|�ǵ�L��~�v �>Ĉ�E��^����P���6Њe_S<���@�JK7л�>J�����r�	�plk<��L��"�Z�k�a��h��������ݔ�1������ୁ������v2V� }�<� ��y�E�Ƃ$;H</�{8�%���0�b?��1��)���� &;F�%��*#��L��DD)<��(4rd;O(h3�Aa��]��c��㑘���a�d�v E>�z�J�HE��&��7n�rD���C&<�z�N�(�x�����|ҢD
6b��kp,j���+�p�1��9�}�)]����B�!��E��cA�� :�J�CY�kd�(��nW��1.���"�4�6��5|ݧq��G��k�2x�Q�V_���߲ʋ�&a��	m� �#x?�t��P�����~���?L7�����Q�I(Բn�&zw�'\��4����O��;x��V�G; ~�?�8�O�X���� _{��B�SO=œOvm22Q��Ȯ�>F�$�ɵtZ�Q{�^` Zl��Q�M]�������N���0��er�f'FTD}��w~>����4�u0?�s�[ ��믳���_b��/�g���}�a�~��/~� Bd����K�&��v�(ϔ�=� 8j�6�#����H��b��b�^����P"�����JZ0b�TVM.�J���y~���p+J����g��;{�%R<�.��5�,��GqE����x�]�Г���c�1 S��w��߲����;���`3�ْ��)�.���	��B&���̚� &2���|:_=G�(��|/m�\F>���&����B0ОV�*�y|F�*�컌�?}���&��ښ��<s�L�P�\QO^�LLq)6��	��l��0�Ђ�r����x��y�B mF7,$�uY��#*Z��a�9��LP�"`�äǳ~���gM���y�~�I�&�_D��,���]`����{Pp.�{�M��rr,vx6��xθ&+ v�9�ոq��Ya��������B�+�'��Xu���h��)%�{1���t��jN�fQ2UG�L�'�"�7��OI��ӀA#�������@�s�@6�r?��@�讶>�M<v��s�����D���:N	���j�Yz`ZI�_C�ʋ��>lԁU�vݒ�!��354���y.@9��|�h����w)���D˗~�Y=M�Q���Z���U������k��b1(�8���j�hъ�m}��7�A�`Q���1�-0��Ȑ�K.I�'�Z�,��t(��Ď��������f`��O~����#�0��?b ���3�h x}�_Z!*���\W�S*Z�Î�B�Wp���N`� 9�v�L���n�İ8��x1DPǊh��B9��7�a����]w/��=��=�=�-���P�K�����1���$vK$�h��h"�t�㬷�t��`�R��]8���A���ߟg�tFb7esB�8�9��͝�믲3���z&;  �k�uA0E�[l��ؤ�z�����'m��w�2�]�a�.�������$��t�]u:(� �3�Mhcp	e��j�	Z�b1��[N>�E~o��Q���'��|;���TFY���Ę�4�?s��=�@h��U� S��16���x�@� 8A�������>~�\�VB��K/����cq.���(�@��Y���������_.��_q��)������}�g����TԮh�h@���{���
��BH�,B(����X�d�õ�;Eܐ+�`��n �� �yj�̺�)�@�����Z�\�?���v�x��<i,E�8�c�R�&�׿.gWϣ�:���	�n��~C1�_�{����>����_BpAD��E3�>�3ĉ��XY�Equ��
�~2g��'2��9|�%G�\�	�E��#����%�.=�K��m�����Ȁ6�����	��@�d���b$h��o(T�|��f���]!���\����y�C����O$�5�N %�֚iDO#H�4*�q�k;���KJ� $�;$�B�t�E�@��?!�4=?��#�W>��w��~;����?�1�eq�<�{�w HaW�����ڴi������T���x ��1�(&LH{��>�"�	�h<�	8���L9�98��-�]���s.B.�+D���u`�s�y���E�w4���!�0vM�:�,� ���
�t���	\u���'R4nq�^s����#�3(�?�r��������8�]z]��y���ϐaQ:uW�F4�p�iO�BU�d�}t#��ً6���� ����x��; '~YY~��;�` ��Zj�o�����27    IDAT�(���ƊFԾC7Z_���.+��0"|���߷O۝�u�t�xa ��I18
� @��M��c)�iUF�����uA�����y��ǩg�^�9#�hZ�׿���TPX��x�hh��^�S���c�� ȣ��,V��@����5cG��K ��\�7���6j�Е��5���of�4Y�s�-C�c�wh��E`����i��c��;�B"FmQ��ZN�;~��zVO��f���NЏLJ�$bI�s�.��#�Q )C��<^������b0�/]�2c//ڤ�� �sYGd|:G����~N�aQ��g??��mP�o����P=bm��
t�1�g癑�Y���89'�^U�ro�l����-j�b�0����!�9H��Q�<������˧X"ɉ��O={(͂�����Ř�P
�/솤��h�H�'5@р�����c� ��9@������y�^��c���`���7���� p�\�]Py�߇~�;�@
P�1c�a! �ʽ8��&�馛ҁ� g|�Pa�B�kKIP^Ai�3��#�7d�G���>��)Y$|C6�},hX\�N�+�K���E��}�$^�I�w�﹂��硔!���R��ԑ��d��~��?Ծ]g6�r��]��J��rTSU���s�EC�|�wI:8Ѿ�0"�� �3[�n�'��􀓟�l�d��X(L(�x�`� `�K�-�X�w�q�_�^�8�'&�cnJ�ʕ�i�ܷ�&���~���~;�Y=��mՒϛ��%܏z�(TG��Z/�Ȑ�H�J�ᢿ�cE;�/���>c��!T�ѷX�la=x�Hv�D�\ �C�@Rn�H������q<�����������<�'�P��*<_Q>����Ba1B;�o_\[E�p/����!��RAN�y�� Ա�by�[�v�W_}�89_vI�����F��kz'����sp��D-u��P���k)�qv[D�#�-�z"���ǞH�����s����<~P�w���ڎ�$��9��f��3;�Ocm�!�9�W��u�7I�늑�@��ud�\=ۮ�C��l�d[��~�cF��ɇM��p��l��2�!�xSL	��N��|ݗW�� b��DRɫ�k�Sgٲo��l5�=d%c�1*H�={��\]A�|�5UVE8�F���Ѐ��Ͽ�k����q � ��N:��W=�I4T�%:�b��X4` �5j11ax=�i���L�`��w5vH&���ջ7�
 ��~���.���i��;���ޡEc\Q����y�B������d`�Q]����?��ϋk'vH���(hY���C&���}�;p�0�"�0��XH$L��+�
	@�	H�*�7�<�&����)i�q��.�\V�*e/+�ѣ�҄	�ϓ�?�����~�~k�}ߗtB����� #�ҝaT@@ �E��8��1&�0Bt=���â��d�I��{-�W�V뭻��|���[��Mխ�y[��=�Ou������<���<�͟��T��FƊ6o�b�����X���I2�����=wr"�ց7Y���D,��zW���;�|���^�}_(��yԺ{{�g$Pd(��e�d�+�V�#&)zF<�����k^�j��h��3aae��3�Kֈ��8R鏍��:`���W���F(�`<=�i~29��F��UO�!T�x�N�d�h�\���(|3��Z�r��{�x��6R�K:���z�+(�E���qu���(a��r84�g���\t��y`>_�!��0G6Z�={\�%��G�eB���#�g������B���8�	��^�{�ġ��ݻ����QQ�0i���c��*<'J��SJ
�;4yNA�%��,�Q�<��r���;&B=�p�"dyw| r�J��u���p��5�o �չ��g�^�5�������`==��÷^�͛�{y�L��Ț�綶�V��P�YG�l���W�x��{9���fQ�4{
�~�w��<31/�(>Y��}2���ԟ�w��VB�5�f�:W*�-[�,�xa��T��*���l�����s{)�R���)�q3�f�@,�f������wO��'">���k�m"���m[��*L����X�`�KkU�c�a6/�	�S,�ȨdQ=���D�;^�[�z�N��ju��Y�~��^-Z�����y�sx����6:V�F�bfk׭��+����]ҙM��I�}��#"'\�C?���f2��į����#�F��ɣ�C���@D4��v]�M�0�c����;~��qo�q��C�&@
 ��ً�Z@])E�KX�S�XZ��}Շ�"�uP���(�1��@����n��5{�!͟5��A�4Ԑ�p3���<�G���z���|&a��y۹�^�-�(Y:Y��n��Z��iu�9���q��24Hi�X!����Ü������uA�l,s�k��f�w(a�;�B�e��((���n��;za�cHpO��:���6�4��������mOJ�6��ͥ�^��/���0]3%h�yX�t�z�+��>�D�N�:a<�]ג\���m���U��\�ȑv7á&��DGH��h��Ֆ����p|��Oʢ������n;3�P��\�;��2���}���6:ְF*��TճQ'R�Ǘ�T�̉F�ɘ�zPYߠq�b��`s6������Fи�����/|�A�Z��U>�s�\���ż��������)@���8v�r]���'��7�r�SWh��L����G�#�'a҇
QE�P*�wı�D;()KB�{f�S��¢�^��L�?Z+q�X�X���c�<����>���͋��7_w��_��V�^i54Vr*u�ow�g����~���y���˦)�@?�e��{������b��ɢ��p�ʅ!��S��#���ظ��x�����v�?|�P~��2Q���?�8͙�e�LچG��g����M��K��ƍW��;<�R��U��̳OM�8	:l��z�>�5���w*�_�4k��K읿�v��l�T�a}G{o�J�d�Lڵ���CL[�i�������y\ D� �4
�cҵQ �"I����w���hf����<9筷�;u�ی��H���;`8���q`�[�Ɩ/���|�����7��K^k��y]�	�Xiˊ�bnЖѬ���7�D�G;&��_ו������	�����?����^����-�ͺ����l��:d��r\�[
�h�0��A(.c�x@|�3���'����J
��p��1�x������c	��@���IL�
�M���� ?�O�u�[V��T3���<q�>���5sI%�Z��nW��F/�ݺuvͳ��|�l���dl%��C�8ξ��x~���?��I����eng��f�XC�x�T@ɲc~8�d�ŋ8M{��I{��'m�L��ǜV�g۬X�x�E�����l��%�\����V�Xa�Q�X���i�={�xhh�����dO|��׿��v�O]���~;u�=�k�ϟ�S'�˲�H�ldp���Z笥����c�S�cO��dN���N1�_~4�OZ���:�)�3���#g-�L[&�a==��U��86��&������ݏ-�Ϙ@��1�R��B�㌖̢��������LlEca��b9��7{��; �X�YE-���͋�G��x�?�2�gh�>�`��gº����7���;o������ODٽ�i�7k�����)18�y^����ONe'#9�6 �� �!G�
����B�`)�
�F� ��/��K��M��ۮ�-�iX�D+G�ի7ؚ��Xjxm�l6�a�����yFm���(l�&Nw��F�}"m��G졇�^����J@맪't��uyn�
�U�kTG��w�����J�UR�V-��[�a6^(��c�v����7���$��_��_��u�Ȣf�'.�v�����/6��O|���=�������&����Ä��}���|�b�U��o��/m붫lt����?�ٰ,5AJ劝<~ʆF+6p�lo��o�9@�Z99O�c�������R�?��Y�<f�d�Μ9b�=k��l��Y��?mc�����������㣈*7���`��%rg��s P6'��E3f�J�D��QCu�K��ht<�?�g���#��2��ٖ�[=�h�O�s��#��ޫp�2��١c�����J�'|O��BOhМ�c�	*JH�� @IF���}�"@H�C  ����]@(@��	T��8��|��O*Y��������K�Imݚ�m���,���*�`=_B8�;:]��5�8|Q* ��z�(��o}���X;U�|G()��k��<��J���=k�ʈ5�e�;�g��H,sK2�fǏ��b�aǎ�[��N۾�j��=��<H�G��d�ό�[���������J��{����ۿ�V�n�j�?�h�]���"���b1r �r����<6`��,;|d�6l��)Z%� ڀI��Y3�ACCӜULG��^�÷2^���\�a=={���V#q(�m��� �i�B�2�>�l��e�F�9��h�܌;>8ru�b���,B�(@���d�Q=�lp�)�+ |��;��/��"��=�:B�G����@�a]P3�?4�# �5Ƚ h-B1�.��8�cD9�
e��\�*�rh�q�����p�N���`9p}�'h�XXD�`A�(�(i��fM��B����i��E�D����\�m�Ԯ޵���%��m�u�Zd�_q�Y��J���HeL��'�X�Fl|�>���@1����o���Zd��Ԕ"� _!����c8~h�����l�ڥN=��+ǭ���}
�Z���=쾉ѱ��Z�����wXG�l;yj��z��S��[v�ghx�C�4Қ�+�W?�^/��ݳ���7��y�c�{�4N(5M�mhpغ�{�����c[�&�I�X���h�T=#��DLl68q�ԅ<�ٜ���p���IT=sq�8lgN���[+�[ �筯�k�����sV_ �_�3o��4'8{���Q�)�q%�B�=�*����P. ��������誉
�g� ��C�q�j�ε8O�;�& .JJ�E�9�/�%�&��r�u��T�kI �x�St���C�����uT��5۸����|3��KY�e\�#
�$,a�PO�8��������_*[.�r�/��յҮܴ�2�v��	�C@5��8~|rQ����sv�0A�1��94|�֔2���r�X "ð��������|�6o�`����w����b���B�n�=w�2��v��/7�S�|�
��7R����۩��x����u�݃�C�>��=�6�j����T�f���}��u����^�����6>Vp��d�l���9r�R�Y����bӎ	�gS�� W����H�4�8�S�Ntc�l�yq����D�j'���=�X�FB���Ȓ = ���z���J���X�("�y15-�8z��[�x�d2���_߻�4Τ�,��TV�����k�������Щ�s���y�����M��Rք�		��1���ֈ�wx|�<�YϦ���u�q�[���Tb�����*߅��`_�g:���/Xow�����l��Wx��<�u������k�o���h�r۵�Z��Ky�Wwx{;Ԇ�������D� ������U�ư�H�D��̄�B��88�}��_�(�9sf��C�}L�wTm߾nK����Q+V������jG�#�K�qԺ����En���}�|bhh�7��=&���������w��_����~�N8}�J�b�O��P,ّ��66^���5��ҫܳ���I6�q��MQl/�+���(,���*��'~�^�h��>���O=lgΞ�������:M�H[6�n}GO۷�����,��l���d�ǛX\<�o3� (�T���&i��p	����څ]\"A�^��N�y�ֵqB�-v�K�I�&���h�uX��.V�tr��}	E�85F�v���,l���8��^=ח�YA�r��zg:p��y���m�%�b���'�k���C͈���ވ���uA���n	+Z�Z�(�T��͌U�)�5�~��W[��o�6+�	���x\����#�4�^4���}L�oYc8�J×D>�|'�D�#�����)����b��-����?y̪��[��2/�O&�e�N���K���?d��s���1�����+�_�p��fjI����gQΞ�i�|��l��%�ޖ���_�+�Z�6�_L?�;��Œ�����Ƭ�t����w�㌍I�6&E����LD �S�� ���jT�W+��h�,sm�<qB�9`'Ou��\)xUO�Rx/��}z�>i��,7:�f�r��?tBJR���M���P|����Pb!�zC�V@h;��&�^Cm\�ǉ+�Ix~��f�s��4��u�P#��s����9�/IJ���P�,�����	�PP��-�f�L�j(�4�\;l��K��b��Y�{����3~��8�{����|.e�zɮ�b��ܹ�s`���wȵ�{M���k	[�z�U=�&�}/��I|��>g��/����;��N{�k~ƅyDt1O�����N��O��r�>��}�ha��S	;5pʊ�1�1� �z����q������7~�k](}��G=˻T�|�/��$���w����Ї'���j%�F�[n�����6V�F�h���sV��G!X4s��e��6tn�N��5Kvٛ�����<B�T��E ȓ~Ы�
�:�Y({���I$B�	gQ���*�P��>Lzil�Ν;c�:����Y:8�̒�W��И������k����k�y�8�E�}BS?����� �ٔ5GY��k~*�����E�7�����e�:�����t�/KA>	���-�
QNa$����)ԶC�Z,�@W���JX{du�,�4���JP7[*/U�!�/��kVZ�&�?��7��O9�R�9]Y�;���uG�xT�����Ȗ�x�t�KĹ�X |::���@�D��������O��!��R����������ر�����;2|�
�v�d���7Jʹ��:�y�IK����s{�E�?�V[�d������w����po�
b�^�ɝ�n�����M	���Ă^�|���]�b�ͷbaԆG��#�|����D#2)�eʽ���c��̳k����L2�rl Ջ�!�VzQ�S<p�lZ8B��r�h���6�&����5��g��=K'1�Փ��|QS�0�k��B�H�Y�v�z3��	���"!.�� ���7���4�f�#&ː��<iѡ�>ḇ�G ;-���}�Ly����.��9�C/C�<�eB���Ofq�<�q�Ӹ���BJ(����T�<%��f�n�g�Q�����-�({�Wi|��u5�Q�e"��b�b�sl��^�'s���p$����V-����)��p�b1�Z���C6:%�(#��(!�����[�*6p��>t�N�������6K4�^_��Jf슍[l��U^���@�,�p�M6v�Fc��h�x��TEB\�u�ַ���Fm��.;sf���N�BR�}�Nۺ}�D��K�B���u�?� p|�m���P/��<0�	�ęL($Rǽ�b*��'�}�8���Þ^�j�ly��b��6^�������M ��������{��Es�����oH?4[�=�/� i�D�6-�?3QP:Oc��!@���|�eYH��y�V��]�#��� Y�u��K��*,�&�3�4����v+������m����L����E�H@�X����,YBmh��F��XH�@�.��a����z�T��W�	��I�ܰ�J��[�yKPJ�����w�    IDATa�1�>0p�>��>g�Ҹ+R�Qf�*�K�w%��P���	�ݳ�+�
֖�X__�=���=4���âF�+V���o���̙��B�9��E9tz��gF��n������_�J�WU�Z��Y,�{ӊ��Fn���I;E�0o�Y���p����=���Q�(&���:���P%,TZ�7����T��@�ؖ���5m6ɲ 8@ǿ�~�N��X��=q{:�p���{���=f�c��f�^%��[�bu$$�+�x�>���GH��+c�����;�R���m�N%<D{|��K���t/Γ�PXg���<��s��9�<r�N��J
�yo�y�B���C��g���ZD )�?�~B�*O�
?�'�����][�P��7P��J�D��U��j�T#�?����Ջ�}�e��͖�G�I���w(������1��"�oo���>h�����y�����w� ����16�C�w�hb?��
7V�U��`���J�IgG�G���%'%0%�����xN�9h�o~���v,��%�Qѹ�>3�o�s���{%�D����.�ȭ[7{���~����{z�%HĿ>���.��nB�S-5�&,�E� `A�!J�Ϳ{��y�E�ڏ��T~tޟ�rq@�U���,۾��@�/�z�liZ?&���s��i���R�膜7���K�)�-.nIg9 
9cƀM�u���D?1��Y�*Q�xJ �2��/ R�fb��p"��P�G`c�q<�AT�^c����9��p׆� #ƞg&v���]�~d��X(�D�l5�x�,lz	M6� �g�W�%����[��{�X��D�����pMţ��Y��	���?W���M%
��g,�G�J��%ͼqnX�q$�AIz/]������	O�"ڇz��,А�y^}�&+Ǽ��$v5��'i�5{�]�e�G Q�n^hހ?-�3������w���ٟ?��M���\@��G���}����Ԍ��E����[}	%oԫ�k˻J��7�I%��D}��oG�qw�tTl���,����i��1������+lێ�v�����Ʉ�g�r`ч�t���A�%ٚ$uQ3���L���OD��6��#����[5s����#�m�T��k%��F-���B Q���}}�v���c�굤�]�>���{�.�CI[�j1�� �f �qz!`�v�V$)������a���G13	U�Yuo(�FF%�qŜ�: !ay��l<
�~+͘��l	��������͍�M���4�H ��zTڤ\��}�A�l\(��F.�$�OB��|��'�G�Y�Ō�Z6�.܃�PuX�EX�=nٲş�h
"@�*V$�+�'������Qh��'�źe�B?��Bk�8� Y`<Ϗ��5�j��U�P�0�{'�����&�.��	���Q=���m��N����^�皫7��)ژNd�TnX�m���3w�OC��:��6��j�Q����g����w�����n��V��#ܓcM�?B����߉R�>q�w���Q�Q@j'��")���ɧ��y@�Jd��]��'��L�󟺼CӨi@e�+CVC�c1���dܵxMJ=������I�' P��?�A��{|)S� �0Z�����j���9}�z?g�҈�57sm]v��xTۇ�΀������3/ry�K���j	���Q@���#��	�c��ËEŘQs���%@�	� 4(�����E�y��G�MŘ�`G���G  Ҙ�gxX
�Q����� U�m�|��ا?�ihr4e">���fF � P9���F+$������^]��C  Y�J�`� ̈�WD�.��@E��]��A�I,�Y#�1`iV����r8l��y#f��C�I�����Ġ&e#�;�G�ERm���<�04ɅX-���� ��$�"��*��9����g��zz[6ٰjm̶m��v��̊��FK-a�L���Zn�6l��IZ��Jw�jO�?<;�V�
��}�3 P1o{���C�kpg<QX(�G�&(�ЂcND)�*7�NtR@O�'�1�¨�h��o�u�g���?�#Gd���Z��u՛9_E�4K_-��-@`�g�e��� h��[����W�j�d]�.��������iTk^ҹ��ɉ�nQ3�FT������.3� '�ECcs��Y��� �G?�Q{�k^��-��L�� F�B[D@0/l@�z��Z�	Z�� 	@��Jm ��4rd����c4��kM�b�U���<� �l� �(�v-.B:g>@(����;k�͏@C�N�0@���Z@�G���'
�!T~4��ތ-��&H��d]!����ð`X�|�*���I_c��cҌ	sûBePH��5<7�KDy��"4��v�!�0@h�>܏�X�|Tj�#'���J:������@TϿ��r)�re�vn�ܶo��C����<.���XǬ�6>^�j\ٓ`	�ѕ�j9�ԫ^6����
���}�{<��g�b	a��֩�
�KM	X�5s�5��q�~���w�5�x�}Z,�j���XͿeU�x�B���P (��9�Z1�!'�̿q�����j���aΫQ�%�ܻ�����e��O����Nؓ������rVk�����#66vk��bY�����{�}������VҏLd�l��y�&
�r���D��� � ���1��$�Q�8x�cs"\��;�U?y>,1�h�9�ȓ���Ei�*;V����$n\��h� *-3P�� k �x���������]w�����@�g=�BQ	"@��L�6M�i����]ԑ�5� f���tPj\���E�	���L l�������a�b��bC��@�1N���xƇ���ȉ�����'̎n�W�6О]�$�����L\�?�ߊ����k��+��}�Wk�^j+�\i�:%*���4�N����LD�`&�t�A<V(x�^��GuPذ:��+S�RZ{�#��X(B4��/֏�����G2�5�[v�~Q�\����hIi�k���P�H�7��\
�G��;�1�, ���%��l��ג�M�^AC�ٹ���'�F�>�ԸOؑ�1��MN3��zRҙ���3�p����d��w��0XGP2l*U�d�Uvm ��PѪ��DB�;>|  ;�8�0�k3)���C@��riV�g��M-M�gCp��w�s�� �?��s"��]3��n���~Ο��������D���Y�\��P\��<��E�@��z��"� ��yg���̀���JQG_,,31��5�c�b�7��1�Z���`e�<ļ3�h�X#<��1Y9��J�\ɩ�B���������|�T;�k�F۾�rK����9��z�[��*�6�V�'�A��Z�����#~�<�b���r�|�9ғ���wG�S_|ƞ�fܨ.���|�~��0�K�-�I��!� ��hi����o1N����wF�����#��T!�#�r���Q6���ߘI�\hQ*��h��X
��h���k��7,�6;kǎ����yR�s����3�?�����������F� � ��)9 d��!�D�������C�x @�#xo��c��E�b̠'�ș b +� ;ԉ����� XC�\_�	�q�H�h68���������@��9~�"���t܃ka)��o�[����g�Fk�Fh��:2�� �j��
Nj��x���NW�AG��}�N�O�ϸpm			F���X.�(��@���c2�|x&(N,+Q��������&�d*Z�����q��1���*�^<����F�*6�R[�f�͞���;$29KT�zD�e,��ɦ]������>_�zT���c��T�9U�g�{	נhq�a��K�F0�\Kʢ"�Z�����n���}n�whh�=Sq�tih��Zf��t�Ĥ9M5��|Y ���hB�)'����A��7��ꓨZ�6j��!;s昝8�cV�!�_	�Kz��Ѩ���>4��G������@�KfY; �$�V\04`�JX�M7��9�GÇfPC�8�~E��^6��0�8�c�9�s�����8D���<#߳�)ԇ6�?�v��X�Zͩ�	x�ݰj��p�h�8����K�X��@ A�`=�}�4d=���7�e�@s�R �yg�1��yXT�3�$~���&4 ŸBc��2�9��	�*����!|��4R�C� �emx�z��~48q����2�p✃pVn��k̉O�S���9��Ba7���{���Q+�V����d�ƸY��c�,a��$;q��<���ͷy�;��h�T����;�z�h���P*<4�ֻ��Q�G�:o�@	;�£C�AX���J9l43W�e����{*�,���w�Tܿ��Pp��C�˹����5YD���s4$L~�^���0KT���G�T�eSu��j�&���NB=�����oT�?k��<� ������4PQ5
d18E����� Z'�1c�E�3�aB�) 8R����	x"Դ]4���
d���V���������w<�V�/4�k��b�p=��`m�vۻ��?BI B�{Q����Hy�6c�?�*�8[�l�J��G0����;����F���?A�T���gM3X<�/��cqM���r,ϧh"�Hh�r�ù�0h$�3��
���'��O3��[OOTҹn�y�Z����I��`Z&=�GJ6g�����a)��I���l��g\	#��λ��9ͷS!7:��yY�
"�~������؇�������l���-Xxیl�8�K�ntw�0�q�prB�j�2Y^2��[��8�l<b���h�o�bO?y�x�?qι4�a�nƶ��0���o����ڻl�P����g)�����S	.Z�DHP�Q22��R�o���3����^�"���dI�����cj-M��C�h��+sqmy9�B�D@������~���uq�P*PC�,��D!�y��XD� ����=Ѥ�%ᫌ�Ve�� �;��b�f�xVU��$r=��wFH��ܛkb0g֢��/���a�w#��5˹ⶹ&τ��傠��X��"��S!C���/њ��D�Oe��/Xo�a��?:v֮�z���S�l�0�;�L֪��n�:V�,���WY*M[Ժ��qͭ{�{��G�c��Oi��eh���B!�5�R�C�����R_g�
��֘07��ߕ��
[�y+����U`�s��ܥ}6[�'��,*�k��Z��1���N����A� �w����W-Q/��fuം�,�b%K1��ځ���Ǟ����'}���r����b5s�F�C�$�Yc	8C�����@���Q�ތ!�E�	�7��ax�"M�0И���$ņ|� ж�x�T�.�A̛�6�^f;@Z#<a|j̃���%�Z� �ϵe١y�
�û���������]є��.PK\ޝwCx�[ ��&?m+�֋�5�D�qo�K�1�r@h��:NYuSh��W�.�$j�ga�3P]�{��	�����Ԯ����=�MĚ�y�5� Z�w�*��^�vݼ�&8��+⪞�"9|)��qGj���M�m��+,��z�o�ޒtK���Za�dU/�\�|[�;~=�2���pl�+|��&ٓ<���\�Q�F�	�sQcr��]�5\g���p�$E�_�F�Z���,\����җ��������i��3�,X����Z�)TO&1�b�i*�xX��X��o�y�%幷��l��Bi6�j���h��IFo٪%
WQ�6�`_�elp�`�D�ʕ�,q�˗-�����0�a.tލ�6?!��s -�b��@	`@q��Frt�'����� T�7 e�����+�G<`�#�EH	\4�2�����hL9^��O���1�z�C[���%�U���yމw D�l~�#�����>Pp�D��`�6M�)`������P.��揟 ��Z�̬]�%|%aƅq@�p<�
M�{a����0��<B�s�P�^�R���A�u�_~Q'-@��\<�g�
/�|��D��Mٓ��kE��H��Ymf����)����@�'V�&��HY���\�͊�(@�8>�}F%�P�%ӕ����(2֒
���Pȅ�(�kM��0��f�*��Y����o��o�����ӄzJ"��*�]��f`s�  �]Z�jvȡ�w �4���S�!�P�tp�:F�)a�`���CV),�m�yu�(EͿTI�h�j����3:-_F���.nw9
%д	xW���`C! T�5 ��ln~'�@�)��#��i�r�|4t�08�*<6�~� x.�A~��&����>D�i��W+B-\�7�E�p}�(izh��MJ�뉱A;�U�F�O<�:�j�+34
�B!��/��%�9Z������� 0��DQpO��\0'�cM2����X�#Qb��S~"�p8�ySY
���r�<>#�V Z��h.�d� �~X4��XOO�u�wX�4b�d��U�4<J[��h���g�Ξ��6n�f	�zE���1��eU/��"n�駟}��|ܰڇg�0�����1d����h3�Z�̍���a����1dO�\�l�߳珇�o���+�����ĝ�Q�d^n�^���t%"�́F��l��
ȧ�Ρ���-\2��*ɋ�'��������Z��Z�D լAU�l����g��R#�n�/Yk+�/���HR��q�Ffч�Ei��5#�_��4om
EN��F����Fi�:�ߡ(�#E\pOi[�V�����

-/��d��y|�dѦ���ϵ���s�4QMat����QD��$�Bk��d���T�A��,S���hL�!ϫ,w���3+��Q��9��q_�%��k��Ƶ5��;O�o.�����cL�8�S���s˹�(چu���K�X�:�e��(y��i��;��x�n�V�}��N_�"h�h|3n�}�'#|h4\@Wc+k�C��;�
�C9\�1W=)�%�f�0D`C���A("4�(7~�20�OD{
���Ok���f0����%����:�� *�y4=8LņK L�
56�xa��{�c!���I&jv��S6����esIKԫ��ʣ-:���}灇md���x������5��bT�x்.��ؠŰ��=���yKi�l,�IZNH�79w%�Gi�y���X���ϩ�' �Uǵ��#%ABBڜ�Eq�l��tM"kI� DJ�~���7O���Z���9�g���y<oi��IWֹ�+t�A�r@r��Y'��X1ךC�'Q������ʟZ�Mt��:]�l&a�ڸ��v��tnT"���m�7��-�=�����:w�9��Yq�lt�i�Ko��;~�-���7�4AI���� 1���"k�c�
&V"V��=QG�&(�'(B�>�Kx%`*v�e�o��3	�+76��8��Xf��&4�"M�c�˄�z��8��H��{Q"'ؼd�NI�$��w�#6<|��U4\VQ�p����a����~�
cKg��J8��{��b���N�"�i�r�3C8��j৸T��j�(|�kl�fB�I�� �����p=6����k���mq���G�&��E �@��8_Z��$��>�X��:N�������B@E��}��r_{�IK0!Ƞĸ�4x����(���}=C(�$����$���CKq* �{Pҹ^����aˤ���!�r�z۹�*K6"��)�\�P��l��e�e�.+V�6,��{�&���F�-�?���>h���֬��N�=e������C �J�#c�>Ƿ���^�Z��QLQ4�����/�����>��>�B�>7���v㍯�&<I)�aw>���޼����_h[�l��wy��5�IDy`�� e*����A��c( �*ԓ�t�3v��a;}����/    IDATU�c���(���\~����?e�Σ�Б)�&��K�{}.V��(i���%8F��%zi�i��t!�0�3��K�4���e���I[�!(�u�*�%���s�kB�c�f,����OBCt����9*�gܸ�'�{*��"ǤK��K )�M�U�c��)�� ��Ѹs=	EJ5BY`�B~ 	E�I��&�?/ ������D�oV�M�а7Z&E�fT\.��]�,�d�lպKl���f��&b��'
�������OM�d(�K��d,�ې�Cd��Y��ɾｷ[[[��mY/�|��q{�{߷����o`Ū��;���a�t���Pw�����o�/h�/�����S��K�w���p�l�D�������Ν0h��� �U��⥫�k^i��Q�)�q�L��~E���ӂ���Q{<9�ظ�>��V��&�����f�L�Ϟ�Ç��b��k�C�g+9v���S���;ԓI^5����o^��¢;H��Zn��n|��@Z&?�'p�w�G�d�:�j����- ����F`���l��d�9N���Ӑ��=��7�D\O�o��hQ$�^xvmx	{i�>F��k~�ֈ�AE�	h$T[�~j���� ��.�z&���%�{zڧT�m[/��;6y���r�b�d�.{�.�5w�e3m��ztl�#���z�j5��l�C���Oz�s�LFY�a���5�ߎ+B]�Xw�2BUٕ+�Y�R�Ju�~���l���V��-�H�u��>�.�|�m�~��)A�L�����O#k�g �V��=����F�x	�¼��֭o��
�C66|�N���޽6Vt�ϻ��='�v����+I�;o����q��r�<�f$�[���Ą��O#
ca�
 Ĉ��*�� �Q:e����ؑ笧�+���\&c�|�uw������6�sA& ��F�L�A�����H��}fuF��DE���V�(c#�(cE�	ILQ��W�6E8'@U�i��[�7	ݛ���*��n���s ��Һe��9
r�[�{Y���k&�ώӏ1����y�$넱iV�uC��z���Um�����q�'r���m���M��b�F�/]mk.�ʒ�v+V�^�'�J{/���X�)K�纎2��Iu|�Ɍ;g�KE��z�����{���g���;�����ș�G��{�<�φG�hR��
R���F+���]��M��	+���hѾ�կ{QH��~�VY�/gny��J:k�9O�_�h���i��?��-Y:���<u��e4����ㅪ=�o��������.�p���夝J��-��c��6�8T�>$<v-7w#m�T�����Hة�����,����$g�ݪ��&x~a7�FKs�����'~��S*VX��ЎD��8�\T�����U�� watl������Bg��q�lB2Y	uĤ�C$���$�!JK�ҶC��{`��k���;D�8%�qo���x��Y�8p��O�h�ٯL�� �N�	��O���d.�?Ɓ�2j"ϼ�S�p�a��/O�U�|�R�Nh�����?��zy��;7Z>mV$,�Ҷ᲍�pɥ��tZ�R��D�9���9���s�t2�@Nm'������=���y�X(z	�H��LrY���?�����z�F�O��O���Ҹ;���Kh����6pf�j������b��^����}��H�iB�_�I�t�\�of�aK/�z%��R���'v�+��$M�{�[�i����cG��V����C�e�.O>Bsd�PGF&�f�_��8[4?�<�Wm�B��>��U+	�fR�˖���C���I�T�L۱���f./,��O���0�����O ��fc�H�v-���������C����p�#:I �Xq��0����>e�)����x^�&d]s�� �ʼV�l�"2b���z>6*N8������%�9aA"�W6̝�"	LDl��u��I��Z��#��x���A[�j�+!X'T�Ĺ��#������Ci�G4�L�LK����C3�-�.�]�l�|�zѬZ��K����vX:�?8��Rz��>$|�͒Q ��4��mDh�];=�\�H�#Ɏ5E2�Ah������.��w����_�����C����s>�POc����{�::�ّ��v�ƭ�����^��pw����:u©ח5�Iv�-{��l�X�W<Bf�ʕ�[��[�j��ࡽ��w��j�g�8��&�D=i�#E;q���>=G���;<}���Ԣ�
�(��d����pO��� A{�yal-�z��&��l�'{��@��=s܋Y	Eu�W�OU����1���S�S��r˥���Xp���h9�È�j6象<���pp��.�(�' ��LZ���'��0��"��|
��tE�.��JHK�秢v�`��D5���`�����/x6�9��<6w��-A��P�L��\_���A����~e"�MO$��:�*�#~r�>ƃ���ь�������j�yrc\Փ6�1��s	��kǕv�5��j��UzZ����m��E���T�?�ō[-f#'>%! tJ�D4e5Ŝ��F�&un#󙪬R�Kb�c��.�?5��Wl��ˬ���{�.���3Y2���S,�j��g�-����;u��M�pj���!�
�̥}��d�F�%[�z�}���3�(��O����W_����w�5��d"c�C;v�U*i�>�?Z��o��J��|���J3FC����/�뿣ɲ��rQw��k�^.���3���g���&�!��N�[w�@Tҹ���Z�Z�}�����Lg"39t���+����dI�h�	GlowNt��elr�)�S� L�LS�js��M��B�@��	L������|<;N;@\8s��]Ř�;����u�������Z|8��9�g���|hͷB?�t��Vu=5�x'��8`��6

�$�D� "N���-���pή��*۱s���-���IZ��0Kϲ��V���Kl����9&��F"�0S	s�k4�.ؙk����	س~Y��]��Z�R@�,��s���y���X.��cǎ����HФ�ܡ�G����ђ}��`���V��Mh���
��8c�8NG��,��d�:�������u��/~���~��2;ܽ��Q�=��C�#v��	�V3�w|Զn��5 �^�E#'��@���h������{7'�ςB�g���� ��M�$��lh�%%�g^��z$��������X�Ƒ�nk��ˋ����
� J}�G�$�86�\��X8/��:G�XDu�0�Rܚ���<�� :�%���c<�7?
J�P��&��͇&L������A�����q��=T���/D8V��!U'+�9���ޔ��܇�D$�p9�~Rl�|#����(�-�$�Ph���z��Λ�q�;
��}�9��7�у��
�]�H��
��$jhZڇ�==n��#v��+lێ+�Ny�l5/�l�U�d���]`۶�Z�J�9�T�lg�J���|��]wOXz�e�4��p��)�֨ΊR��l�)|Sp�(}}{��o�/��ʵ.zz��Z�!�����Xɞ}%`����Y���5��5�N��v������T�`����f.�3|�!��-g����ys�X�������֯_i�cC6<�OF�����;f����l�n~ÿuPB�S
�pO@�C��P,V��͌_Gi�L.jD.���E��M�qPKT���'�H�~k�S�d�3}]�E�I�[O7���9�����Y��<_��W-�kw�zʣi�_�-Y��n�G&Q|7��MC���p���h'~2n}��@��]�M!�F�6 ,�	�Bgr�+�J4WsC.�6s#*Fs�d(9�$�(d��z:j���J��C�b�K����8yk���߻��.�8ʹ�����.�}>@��%��`�'�7�}��1��_�mۖKm�+<�'A�;B=3yk��l�P�9�ث^�+)~����~b�� ��wMT��C2( ��)�>�$��K��`�}�"a�(
��=��7��3ms�̲��38m��y���#�ldt��O���ڛ�g^{�7�yv�>/��E,+�e�o�
�U�L��J���M7��n���f��k�#�$h�,K�?[�9WΟ�S�m���������S>�Z`�q�UE8A�
y9���'��aѱ8�j[��U+E�7��P�8bV/Fez)��ى���s�mx��>�锭\�ܖ-_9�����_�� ��r�~�~�ߏŷ|�R���W��Lԯ��"�І� �z~�w~�#��}����&���f�`m�	�6�h� +?Q>h�,|��\���&��1/8e��XlR����1�jnx6Υ.��k hb|$4$,ࢱ��D��I��d��q�a����PH�Ї�}�O�����w�r5xq+%Vx?�k��1�k�߈�Q<7�w�>����V�h�t�๰4�o���PP�;���M�>�a�C�#Ը?����Z
��x�� ʵ'�L�v���lTҙz�����_��.�b�7=�륚�sY+��R���ZmX�FV��Q �RX8��t
�>N�5���N�@7���ظ+����cL3醝���s'm��Y�JH������1��=f#�{ǯ���`����}��}Oa�Lc�-X��/���|�L��9u'�F�J�Zd��Kv���/���6����s��SO��J�FTK"E�� �,�]���;V�dTT���Z�1�p���lf���" �=�7��b8�y�RqI�L1���U\@5j�*{�?B�\%3��,w����96^"d�b��|��X��
�޴���}b�R�ģ~�	���t�Zf��t����h��i�X�� �u����ȣ�� (m@J��!c��� 8����В�3�X���&��y�&>;Pо8_t�TH�iL��9<#�}�K_�,����0f�a9`��� �`��B@vZ.�l��=�Ԧ�	�L	`ʈ`Ma8��J�v��: J�φ�2�D�!�yg������.X���˚�3�Y�Șk��z�|x�3���5��FR��Nh#��yg�@�E��q
�yE��T�a�^��d����d�$�����V�|J2ac�g-�M[��4��z"��(K��-�J�*�/{�$<q��dv��T����xG�Sy:�8S�R�(41�˹0d�iPT��[W{�|�z���(�uKeӖMe�\%���i۸y��[{�c4�_�K�7���Tz��;s�����}ph�]2��xs��HZ%n�<>:�����z{���R������������������a�V��׾�&K��zł����U'���bƹ�4���'N�t�s�� :6��<�q�8M��mu�?q܎�v�?�%��:��L��600l�t���B�
��X��J��:c+�'��;�t$!pQ�����fuL4� \٬$_1ԭ��"d�D��%2�1@�ط�9S(>*��;0�h4"���k<_���ƕ1Ҹ�a��3��x�d��0[��b�)�E�C��*j&`I�c�I`�d/4Hx`@��[h�p�1T�7���������h��8����XB����.�hu�s�?����ܯ",5y8�G��p-|Mh�{� `�����u m�lƁ�&8l� jd4Z�\�5�����>��D�0F��%P憹b-  ����IP������V}��k�9s;�R������V'E��t�=�6o�f�k�v�Xs)��	�60?�G>�)�(�x�b����%HY袁yO�x�޵Ò����{�g�'�ǎۙsg<�c��Ev٥���l��n��Dʾ�������}��E=^�IF`:����|AΛ=+���|s]w�5�������>�4�����uk-QoX�3~�644�?4�o��f��h�y�r�ı���h"^����ب��	��ھ瞴3T�L�,��Y�R�Q���t��C'�������^��s�-[���5#��Bm������,b�n"�`D''�l��e3�b����Ip��Izcs#h ����3O=�&36r��9��	P#�µxv	�x������2��46-V
�E�/Z4��D�V�GQ�G�]�[�/�����y��Ra�� �x���&ƀ����# T�z�k@��X^��>�4��LX_<'�������1h����'?� @#��C�@� �8�Ʉv��������Zg�c�Ag�8?� gm�[�_��`�P��(@�o|��'�SZE�fj����P��>�4���2|�N�@��֟���x��/Xb7��j#i��:���eg|[<t&���½h�B�19�qd3��#ㄦ��\'�(w�wݾu��!��(<pp�����  W�Zg�]�622f�]�큇h��W~�H�L�3��۪�{�0�h"Ж	�$������WU�^6��ѱ1���v���kAl��,Jܒ��F�q|��؀���������`)@�xDJKͿb��>j���d��5~*�B��l��=���=aC�t����YV����ޭ48����Dҙ��>���'lvx�
`ġ���O�k_�:s���׿�5��W^���F������.n���ccqc(�l,
�b�� ���>�FT�]���VZ/�B�)�/�e�h]���Q��SҘ�8t?~z</c�,nE��,<?�����C <�ll| Dƒ{2�h��?����k ё�aJ��̀P�3�!<?���&c�u��6�;� J����F9��`y�����8Xdj􂠅��:P�Xm����{� ?]�L������"�Zh���t_j_U��^����Y&I^J�Ն%3Y�d�FƊ6{�|���<0�.x(:XfШ�?�K��p_�v�ڭ�[@�yG��S�>���������׽��8j���A��j7�(a�"s�\�H��������w��Q$*�MHw�O��(�\🦍#`Ƅ���h���h�L�Wl�-���Ƥ�_D�@E� �*�M���j`�"�p�hЄ=)a���Xm~�v��ΗҎqJڧbGz���'���4�Q�!w�&��p�){��O��%�;�Z��V�p�GV�T�?�@ |�cI{g��n�J���=������G�,Z;|�-������Zԓ�?1�)��q��c P�u@T%m�t�����"���wm8�ņ��A�0�r��@��.aYO�<��q�D�@�BQ>ʁ�'�O�K�s \z�AK���|���s�m���#��oG��G�=���Z�ǃ����f�l�a��5�X�PwX�� �h���g�0( �\���u�څ�йV�� �=��P�Ϛ�jb,v��I�'��xX>Z��͍����f��;��{�r٤U��z�z۱k�%�eW�Ru =m�ɜG�\�y�ժIKeڼZ�C����G���}��_�E��G>2��b|�g,w���*ժ��,T栽c�]q�+�b^�v��x��G�`V�Ç{���r
S��N�
��gl��t�>��,2@�	Ne��F�*e�1Z8v���j�}#��бǩK��Y���9j "�z�$XR��?Q�BB%�[q����lxp�FGO���i�}(E��s�Ġ}�[߷ᡒ�ۢ"j ��UK]�F�i��cݐ�Ef#-���/~8e�Xo_�or4B4M VM�т�� 6���骫� �	�-	m<�m��;(��h�|�8��8��^e���f���]������N�7�6�W%P��`g�a�+GA�E�T\�(#9|�;�׀��g�~�%�)*��b�������}��|:
c	��Ppli<*�O
��u�������r����sq_���ZQ�@�J���zrT+(��eMqM��g�r��8^TG���O��Zͽ~j>� ��)3|[��v�����
۱sS��e\#�?a]]�mΜ%��5�/Yn�z����?�L�ӗ+��>�G���E@~�w����)J C�bY����)6R��1    IDAT�gfnU�;��f�%B�#b�����K/qg��X��A7��SKD��{ǭWy&/:���?s���;��/Ȓ����'���ظ�e�У�^�s/��p
K)Ւ4���b6�������ܤ~�m��T��tf!Q�`J�oDF_[&�)�=m�O1_'���#>n?�d��H[�T�K.Ygk�E叧4�X�{ m���F�n�3.�0��~�X�[Ex�A�Y�߷ϳzh9,l�� F@���G����E�1D}��|������A�I!P,a�Q	�ph> j�N,5Ȁ�����>����.�ڝ|xfq���tM����a�����W�ʩ-��+?s� exVh�2��zr����"����uO�����&|P�z��»�""�k=N����h}��� <�ƃ}��%�����; ��<�s4��/^Ѥ���h���)+m˖vݵ���;!��x�ƆKw��+�^��;��A���{�tųR܍����r�{��`3� (���r�χ��KOF9@h��e�q~'�8B���3I�����"��C��7�֚d�f.��t�Ʋ4�x�ġ�?��g�b�4C���D9hCiSPd�@5@6/+��s�펅%z�Ο�:U��H#JZ:��.^�D���{��g��+Ke�Xo�I{��ld���Od@�l�b��}����X;:�"!��c����B��[�0�<!nJ�
5}Ox�{Ȇ�����������T�V�-����t�{7PÇ�P����59_�V������\�MO�)`h*��s��
 6�j&XQE����_�U6�m��6��::8Xq,����/��}�����d��<q�>��(×���d�9j�� )�IYq�d�/��V��l�R�uJ_e����q�6I�����]�=Y3�j$0���Q9q4�tsnTc���3��?O��1g�k�{p��-{n�����`���y�����y�'6������U(  ������
����� ��V��  	N��h��4�G�U[.e4j:v�:�Uk�3���}���>j#cD-D%�q��\N8be��Sq����.���=����*m�����݉R�g����N��V�2^i���xL N�WtL�M�gCX�D_ hy �)�ĵp�J���j� /Z8<59��f���¢t\_�S?��'���%�-����Z 2
��jG7�waX_3�s���]iU
�ў1�
��ϛ����q�Į�f�%K%jV+���ˮ���7Z�Ay��[���(�V�|�#8{�O�O�uwT�5��=���DAE&)���Y?-�gk#0�YPJG���r|�N���Kj���{�ǳ��<ON硝�x ��O@��������ln�"�Z/덨�U˦y��uz�z�z/�l�͝�ǎ���<�Hk��zfŲ�����2�3n�ieq�}�t ��C/8��Ǌ��Xw�j���CZd�I���55�ԊQ��6���e��qܪ�W�O4x��AX�i�xm��F���vQ/� @j
�ć�Q�ZΓ6�spO��p�S��X�PS�<�P�#P>|G�?�1 b�1;��$!p��_�z�mW����N^���-���s�c�ev�u[�V-X�Q�J�jK���U�l����6^�z���N�d���8%ӨW�?������#���M�ɨ��9�J� �&-�����?�9�?���5��[&�:U&B0���⣨Y�1��)Z�`�B ��p���BH��o� ַ`c#gll쌝�?aC�#�6�JS5Ǝ�L�?U>�5����eQ�H�M��3�ȑXuax6��lt>ߩ&>�X��H�
Xm(ƀ(�ƈ�_Xn��f;P��G2!�d��A�uE����	��P�#A��ɠ%f��!�SA7q圏��kh�xo板au����;B��@Ӈ7��z��Kr�	Łkആ�x1�J?�B����ի�z�o������`==�Q���]��J۹�
�L:a�j�R�v[��޽Q�\M�jn@����I�әk8�H�'��"��d�b��6�<Z&�|�=�|�%��.�{wk�֙��/!p���:�VB<�ł���'��3)� 4�?_�����R? ��؉���@�Ɔ���G%_R�6;�7`߾��Z�����4�˗��ZםJ��Z �@,*%0�|h�Ӂ/K5R�m�iu>����ب	�H�Nw�l��ę�6���G�����P���gW�>�V�6�=t�J���S��r�</s�ld���Y x�Y�sg<%��.�v�۸/V � �Q��t��O"�_ Z����45p��9y��7�|��X#�s�e�u˥V��{�b�����*ik��U=���*��oo��J������׵�����r�7�H)�\���i�_�������6p���!�4���F�hB#�nr�'�جh�a�n����q��4K�-�"Sr��������8j�Ҙe3˥��]�;�w̱#����S�BUh�+����ΪY��C3BP >��je��8N�p I9V�ĮPs
AZ!��C�C�V��i��DA���y���ID*a ���E�*�F��(,������~;��k����s���������_/�!�}Ё!�F�^����?����ʃ�k�`~�����\��������f��A۵�J���͖JT�FD1�n�u��x�f͚g�]�j-�-��p��{�R�'��:�%I����)�p�7��LE�|&���[S>��(��S8|��帝��A�C�h�>��Xlbi~�z�@��V��^{Ķ��mլK�g��Jy������j%��LZ[{��}��~�)�4)V�I�'��B�Oʣ�������y~�a�TdC�Zn�y*�G �	7�+Q�l�i$����xEIp�q�M�Lo�O<t�4q<����&��$_ׄz�2�Г%#�E� �*�;��է`)�@�yF`p}��*Ĕ��0���r��B	��@l���.8|U�'������s4pﵜ[ӣ��o߶��ch�J8��Ixe�f�����M�Z�Y"�v�8U]��'�G=�{/�]ȘJ�z��T�P$T@��iGd����i�}��}�����00��(�	���&�\0	/c�jz�5e9��kG��d�h��h:m��wl�*�#F��$��g�R6{����B��J�l6��˩'ν0�������J�*��c�㈆�����w�C�1/p��7p� z�(+��8���y*#	���&�Fq�Y(Jl��⚊D�#Y��r$��g�A&6�|���0�H���r�9��W9�0�D������h��=�x��(r-j���h�{?�E�,���Y���,�oV+Y�2�Y�:,��rw��/V�\JX���L�ݪ��er9+�"���~~0j����z�S����d�˼`�[����jg4�O�O&_��f����K��f�vv���8<<��ZWW�'Zș'`�����W�� /i��AܫUy?-{��{�"�4j$$%��5��.�'��L�#3e�j�8Y%���w`���ݿO����
��^@4�v���4v� E,)��r%1�/JbGCb���K���`��wfgg��������~��eؙ!�/��s]{�Ιs��y��������4�dh:wx��܇���K��s��P����9�D���}�)��H֬\�bi�RP�UK��̯Y5V���M-�m��,;P�Z,i�x�^ۇ�<�\32���*cS�L���W��/t"4`��ɣ:�.0���
:=��9��������Z���}F��?�����2|�s %-%_{{���'�oނ��h�bkjn�b�`'QX�����>셖��Z��mJ#`�ʙ��D��~�]1�p�Q����G���?������Xv���ɘ�ke��b:�����%;|�۲y4#:=Ǽ�ϼ���/����E�PE�g}�$�h<<H A�?yF�=z���q��#f���>5/�]�	�36y�Xˤ(�V��Y�,f�B��?�.��f�B3���h���O����G��?~ꖺ�&�!�o~�o��@���������&3]rT���j����cC����Δ�o�׎>f�==~��Jf7π�?|.�?yʤ�x�?=t���f.$q�������
d�-[�£+H�bQ�z�=�ڹB*�&�v��qkۿ����7<2m=��"�H�!,��pp�*� �?8OTI�7}�fC^��}ʶkףv�s���ojL8�{נXʒ�&۹����v;q�ߒ�Fw`�@�3;������q��#N'���E��f�Q:�
N�@[I8�
���
�g���
�7=Ŀ�ᛈ�l����v�RkH�;|I��KY�T�ɓf؆�[��D�56��8�b��e�X���S��)E��:F�i��!AHTAx.o)�''>�/k�3?c�L��!������d>�
�B�f��zh�}��o�B`�ވ����G+�f͂������R{�e/{��$9�6V�y�R�d���8���9,�xZ���X��O</U��%�0d�ǆ�4.��i�z���ݹ���>dU��J��V��KZ:�b:���������[��٩�ٳ��O{J	�����U�S��M�ld���#����B��X�N��u��7aȹ�>Gg�4���RD���5�ym3���c�u�e&��S}�y�_d�
��)��i�4y��=4��t`8�u���J,@��<���=���(�¿r��J����`-#jzz�F���������>�;u*�&�yt�����G+�K:"Mq�^��^��ߴ�&
d嬘�z�*Ijjij�~!�7�_o�c�Y�q�;R�i��z7����&Fm_lJ�aB�9��C� 0�}�$�{��>��������:h��)��oHc�P,Y:�jm{=%ɋ����-��>8|�?R�/B���Ĵ��8�t�OC�ۢQ;Q�����}��Ϲa�7��S��$��F��ty���+�T�ui��5�wcV,e��u�57�؊U�,f��Oo(�G�m�稱��~��?��p�(@�ƴ'e����Om��Paޣ���D}g���%���T �����jժ-\�ȦO�i�M�J7xe�}m쓟�����Y�q�uV�>[�m�����Z�
�8aV������������y;�^{��?��J�R�FsC�]�b��^w����$�P7 T�=��s#D�j�rS㇘a�ˡ����|caRu2Z�-/|ڱJѱ���tٱcv�H��v����Z,D, ��=�e��+���T���s��
#�w`c)5D/����y�_�.~_a�}E��2Z��#�����xN��������>/�y�J+��M'�&mN-=�V��d�w�
eknj�dH�:d�!�1V���GA��د��Z��l��	����G��?�yg�r-��|[6��B~����:w����}���㌍�0�^��ټ�����Ŋ��=�ȣv��
�CB��.�?i��t�m�������xOo�ug��B�Rɸ���/�+.����Az觶{ד�L%,�ΈU���ռ�ґ�ݶh�{�^7�%J�I��ۭ�B곐�T�;������g�d|l��r�$��/@����U*v��k߷ݣH�u���{��6�CcOz�r���>Ϥ��(6>�����ƣ�Ȅ	�|N��Tq���F>/:8j	����C���b�97�g��v��\�_m�<`kW�g7���d�j�l��O�j�nt��n2��3C"��D@!��By�������
�l�r[�q��� ��@�6
UpaB&|���|�j�(��jκ�qő���sߙ�6;r䘭]���ѓ���n��K_��=��9�i_^�u���oV	�ل���}�-[z��
v�}w۬����T�:�a�R�q�%�iJ��;U�W��k��/>��� �$qू#� :,�Ph����8�}Ī)K�O5k�N򪞅b�'�466[[�A�����=A��@�ޣ�����o�z��$y1.�K'�W��;�E4u��te��2�yM�bcC�\�9{�e����h��%���=6X�9�ۜ�X��6oZm�*��kV+Vm��%6k�*+V�V.��Z����ӂ�G�� ���G�b�[�ƌku*�� �3�u!���T�_�?e?8�rΎ����`:;;,I+�xh��Y=|����g-�/����fϙg�x���;�5(���>g��m��zz�����[�O�<���G�q���������9z��zp����w[��#�y$kK��R��Z��7�<�4C�P��B��ҡ�����]��<l$6E�p��覧�l�z��b�͚�v�H������}��W,a�;�����S{��X���i��U��x�Ё�+_��]r�e~ppӺ񢋶�&�l���/�9�a��&�.=CY�r����-�0�c�S���+���˸�r.��Z~*�B�V�a-���/�t4F[y
��U����������*�Aa���>����4�Ud-���I�ɀ��i�pMeG�*(�.c>�x����E!ߌ�M~�9�����-ާ�E)K����՞Pb��
���p�O/���f�b۲e�U�}�L&,^1�>k��Y��*��b���:=s= ��Y苡�B�����2&���y[�]�W�������N$��O'?U��_�����'��&Nh�	�Z��=���Y�6Y6W��;;�RK�ɓ��v����rNM�O�3�x�VXt�G��,�}F�PՒE�?w�]�u���>�����]v�k=R���C����fX2��S������i��q�V������R�'�:��fs���OO������'�����r Y�7kH&,��Y�������;݁��4���uڽ�?d�\���Й����z���ꆍJF�a���osС�O6��m��^@G/V�OMz� ��9P��<(<T�) ��-0侀���h"m|���(�34�@ 
K5v�q+��ļh��V�ͅP�ƨ�`	�A�Q�ƭ�b͇~�<J H��Ґ?�s0^�c� ��:�� ��
�1N֌9�s\�N��t�%��4]���ֽ���u��C���D��*�%�,0"�O�흼���7sQ'���%��X��+ϳ͛WY��o���e?a��]��;y�����/��͵r������~��)g��⋼�<?
g�fCP��৒��g����}������ov�sm⤱�c�ϭR����l�v�9`k�����\���B�x�����=%S=j���Y���>���[���v��U��@�}�߰�/�`�X�����p���Y;r�U*��v�5L96:�ޮ�_�MMo>� @�����}׭��8��u UR*��%gt��J�����}����SGͪ��h0��X۳'8|��g.�����!�s�h(��h'����c��<c�={���;<�B~�֕$�ѺR�BQmz(�I��(xHs�ʀ��F#�� �� �!��Um 	"��Lt�+�O���{�nc0	��J{H *������q�"� �p��B�u��2~=�,�cM�^�F[����?�HT�%��c�\SV��������e�N8��p���u����+��P�!��6�X�p����o�8�4i>��x�ɚ�L�ISfz#u2���N�C��g7̅yt������-1�G��G�O�'���g�+�K�X��ڳ�q{��o�ʕ�l��V۽g��$��Rͪ��=���4���'\���
�U�yٮ={�'����G2Z��Po1X�{�����?�^�ɪ��>�����L}���'��[.�#]�A�G��ѡ��,"�J
�PP��8|��l43q�j���<b�o�`:~f�OX�T�LC4�x���i��費�}����&�T 5�3O�����P�\�4s���6���^�!�P9\�k�6����0c#���)o,�|G7�6�4h��@F�q�'j�*�,��QPR䖛�ޗ9lE*�vQ�d���
n����S��PU�b�    IDAT ƳH;}$@�΅��h.���q�
�|J�������o�;���X��yn�8lֆ=�ƪ����T9������2�%$������{�{G�uGC�����z�۴q��q$��|�X"�%�s��G�<�"�z�,I"g-D��kh��]]��=�Wu@��8;�[@YC�!H�f��e��٥p=����<��~������ĉ���m��KE�R��lޏ��w���2������A�����mFֽ��9��w�?�GkK����&O��η�n�S��Nul��D���T�:1`��d��/��^�җ:xP����o���'u����$�:����k�7��m�ڑ��<h����&;S��//��'�#��,�Y*�|$�D�G�9��I^ݧr�L�X�Z���9�3�|��_���_��_ٛ��&[�|���b��Ǒ��9��	~e/+�M�T4ę�( �
�J���h��p@�4K��z��4z(��c�gS�(W/*Jܺ@?��.!%zHt��*����BF 
�3o�>�����{�y�% ��2�����.�2�c�ŵ٫p�\KN%D͝Nn,��O ���Y@Q?E�ϴF<�z\h=�N�g��O�{�f�qo�N��WY<^�r)��=e�c��/k�c&��/~��*���O�;�D�P�+����i*���Y"�A��F�'��g��|,<�����8��}�~t�]6}�8ki�XGg�ˑ�PW(�~�C��ȱS���o/x���+�\j'Or���/|�N��v��|�V�YL�����&�P�xʶn��^|٥��sº�:�����8y�ʕ�%q+{S���c);~�{���&�_��5N�pҹ��ˁ���~���XhWl2{��A�_u���=Z��r6ƦM�BM��7<C$y��8j�	�$k�JIgw8�c�δ؎���;��;g�t�K��S�'1�#w�Ղ�O�UW]��� @���w���C{��"��j���E]��1����-��0�QJCܺ�n6���Ґ��^`!MYZ��q�9�w�;E��q�v���ʚ�`":F<u��$Ǯ��k���`�~Y%|�W�bQ;r���FAC�X��`3$��0c�,9��ή]�|��@�{I(���[ȱ�Ϩ7��G�,YC�LtMt]~
�7/��:�|:"��×f.O�}��_��Ų���CSC�J�|�y��Y������V/�\)ǩ�˜�7n�;~�~����zg�@߲�?�я:��<+����}h��h�����u���u�ú���l�+������	;��k:�X_o�^�����f�2v���; ��*hρ�(�݈v�I3���׿�Z�Ҿ:�ڮ�OZo�)KRʙ�o޹'i�J�j��󗬶+��!��D�s�{�8�}� ő�/��O��/��n��&w&�Y�!g�{��(�U����W�R�Y:�D2f�b�R�F+Wv�D���5wX[,f��p`f>��>h+��7�!lj����r�']�|�;��!��gy@���A�C[=r9(ꔅ	ˋM�5ѐY>��h�(�A���|>�;c D!�!�9�X�+g��|0���5U���" Y'����Su��S*Ғ�{��)J�uHj͹�"���s-�s͘��s4K5|ѳȂ���]�z���&\�R"��s��PEX���H�p]�IT����v(9o͙�>��Ng�)A��D��(E!���8�-K��J`�4E��.�8�O���~)�L��榘�C�D�O���|�i��U��(�@Ѵ�eZ\�O{�>��+���A�_��Я���(+KJ�g���I<���jլ���i���Y6G���G�Bɚ[-�/{��qc'��������;��A��3ٔf6jU�xh�H]Up��ۅm�9�j�����O~�#;��a�b�-�;ޖ/_a��l�Y�X_߀o��[�V�?8|�q�I����?���]w���x<l��f�\(���G�;�k���Y���T�fU��d��h?GtO�,��д"�$V%���U=�|F�d<�&Z?4����N>�ʳ~�S��tTϏ��\2� �Ќ �K@�"��B`��}��ph�'�y8�&�$� ,�.-|$��0�9��LBp��"hq���c�)��cf��G)cz��\�3�G �<��3���Ҁ&���V}���K^����p/��K#`"K.v�ʘ��ʕ+]��pD������sM9b�����d���5t$��{�;�\��9���5`mn|�y�����x������e�l�B���`�����݊�8|�	��˖0�Eђ���b�X�
Ţ+J�Z�&O�i˖��J~?�%�I���Wc#M[ʮ����u@�'�����W5n	tYV�=B��[�E��ﲥK���wn�n��~;~�;�)�BH�̙sl�ʵ^h2F��Z��o_��/��t��s��!0Z=6�Lu~�u��i�F����Bo�́�����k�X�&L�ds��3/�M$~,�& ��X���ȍh�lG�I�r/�o��o�q*�tp�}v=�����I�Y�R�)B��ԩ�=��V��_f��˂�l��V.#��8��WB	�fӽ�5�sڈ��9�����;�0ǯ�إ_��W�Y8�D(���@���>g�|�+�
 ӵk�:� ��CMH�A�O^UNB�+�xrσ%G����kD�5k�g��0gPvX)j�~�m�����6w��hx$��A�%�C�@C� \\��B����"��p=���q}� ��? ��e O(@+ׄ˿���z���گ9@�RB��<@�#��Bp���[n���F�+���A(�,W, ��A,� ��]����g��,��3��E���������}rMX#� ���`��=4[��ૈ�D�)�oO�2|G���[8o�-]�Ъ%:��=I���R�f3gͷ+.�;W�����)錒�X����=uʱ��y�E���u���/�gy�����\�
�8C	y�k_m��u��\(�Ѯ�v�P�𠱡�.\lc�O򂊍MM��?�/�v�ϕ�h�轢��^�4����$+��~P.��W��!�6��M�ߟ�����������?~Jq�lT6?}aqS1�
�\���_�ʠ�)� ��X`��\|z���_�O<hǺ�[KC�J���ͦ�Ix�۾}�=��G<f�B�C�jη���
����C����׿Ձ�g��׾fO<�sOhan���@q��!����t8�� _��v��)�2�4y@Q��p,�\��ܓ���'�=�y�s� ��.�`ܙ�\�w�֭x �	5B��9����T�y��b�/�uh0ƈ?��lXH 4���S L�}XX '�A���l�F�'���	��!8s�<#τpŢ �����ٯP��9����y�#�*G�o��o�}X։�@�s/�k�6�����,����1�&�N�}Ü�̿���ꂛy欈Fb��'�)����f�G��h��v4���Ϫ��m�ƕN��I_��j�wĬ�e��]�Ɋ%B&���|ɝ��7�C�;��n�[��H�?a�$Wz��ST${�3L�?���Žy�W��J�9a�Xߋ�Jy��Q(S��[=���;��g�5g=��h�6W������ji��0O��!�K���D�������^�>��x*�>��'o;w��~��v����2�i�p�ho�xh��o��MZ �D����}?�
��hh�̑���l���Б���Ү%KŃ�_���j���{~�����=�B E����B��ac��‿�s����::� P|ի^b�=�<�����h� 0g^8$r2����a����G ˈ�Vh�h��6 
��ÆF����%�!�   <րC��"Дo�sO�t@��v�o4~�eВ0P0��� P�V��r`�,��5f�h�h̀>ό���	B >�3�@�4N��5��'�)$F� ��AX"�����Cb1�>�����D�p},&����A�#�{"`���9�^��.�'����#9��� b�y&4c��Dp` h�OΎ"�$ ���;|)�P,���5K<cߪy���Z�a'�P�z���u[,�i�r��u'�' ����?�1����,�ٳ�z�7�6���|�c�R�ϣ\$@�yϿ�.ܼ��iTidM�p��v%�$Mŭ�ʺ�w&!pVW��b�����y�p�O��Or>�is�Nu�9cƌ�C���lX���~Sf�Y��ϡ��&����CE���� ���Pa��4��p�n�R�֒9oP�]���x� �}8�2��,^|�M�>���G��PB[�N���k|�2'X��O��2�(���������{ #a��|̫,$@����3�I��������Ƽ1���
���so��f
�:tȅ��ڱ�rJs]@���1���9�p#���c�q�C�kG���P"$������=� �'����~ m��S��Oh�B����F�h�PiD�(D���[).�`yp=��8q�<��ڡ�h�X8�)��E�@��B8 �/��s!�z���j��=Þ�o�`�Z@X#@x&�-
7)oӦΪG��9ڇ�ΔQ�$����R�Z��W5|l)��B��1c'�KVX2�h��R�Wt���op���|��.(YC����}���d�27��!�."���f���`��R����B��X����ΰ�E���Z<a}�Hk�^g5�_~�����j8�?�$�v�"M<�B!;�~����t�oEˤ��TZ��B��_��_��Dy��C��h�����-�q"z-�x����U=���Wky+�؞}O؉c�,ӀI�������j�,�ޤ�+$y-�3��V��h�?�q�$y�I�1 �}�� D��PCc( Q�Y/Om����������I����Y��]�Ce�2��e�?�C�p� �	x�
#�@c:s���4n@P�|O��1&��[�L�#��z ���@`��h��A	N\�ﲏ?ό Ch�>��2V���%��7�G��X�D�H��3
I�E� <PMF@]{T,4�dyvE�)Z�9�|ȷ�ȗ(��'�s�gB�����{�L�nY����O�����5��zl��e�y�*���Z�jD�4�،����ɳ����C����k�t���y�5��S�7��>*���<ɡ�{�_�A� �a>�'='ק�K�ۛ���!D���+,s�9E���r�����2���=|�]񩞞�7�nB����Oo4B:}����K[?8�нG���f�)'���q���9�8���X@1���5�{���G�R�Ǣ����s���ai	�fh��n��v��S������>ف��b�:�/�&R	����11^LN�����(h�������"��?h/4>Q��h��1�����%=��b�a��
	�o
)0E�ֈ��'�(��Xt��U�d�H�(�C�T+�� `|Ou\��>�Z��\GQR$����r=��M֤"�؛\K�+t�g��*���r�!���e�!D���h�|NJ��#d���?`�gEI��<p-��n���:��b%p�}��i����y����}�+�АIX!�m�/�u�.���_�ڤI��${*=�jP<��;�G��@�<ɋ�?
������8�U	���U���B��u���@���38���8��h>���i���@Q��4�)�&_{��f�������I�����fU̓<�0s��җP1����7eZ���wP�OA�
�xk4A8Mi8�������>��G>2�@h���*�v&��"a)KZ���L�b]'xI�b)�<���?l���'^�ڧR�;(�R��p�����p�vc����b>p�AO *  �Qx
��ϡBbJ����7�����[U�l\��aN�	3~Ɔ���@B���u|�4~w��+|
��;��X�@��*?@Bٰ��W������)M�����ݮ��{K8z_龾A_��q�����T��br�	�
G2t����N��!����G�Gs%��s�̫���{�4����SF5SM!Q�Q�$���[��8^`k�,�t�jTM�C���KmּU��W���d2�)-$t��hL{G0��sS��O����� e_�w�5�Y��`-�|� <j�� �J�=���u���zC�
�J���B)���z�s��f��m�>�����3j�5����^���
~BX.FA������]*�tS�8yN�IT�d� Lp�*(Հ���o�;~0U����UճZ���=Cq7�>5J0c2;z�ö?��� ��2����{?[�D�����/tǫk6�vc�\�y�X4�F�I|���s�� � Z<�,��CX��@ �
�s/zB�%��i�:P�'�4DJ�LS~���e�&d�E�1i_|A��4Ƭ���"��rUn�������wyN�/��Z�l��D�B��A�/E���" x�Q8���e �������J���a˜��+!-Ag���|f(x�<����tV��Z�B�������B��p���S$'g�-�իϳT�j�R�
��-\����_c�J�2���C�Fē�z��Ԩr>��W/G(Z=��,Z��!�'�H�#��u��ϧS��T=��s���)�����M'�<�s��030�'b�$n�
�w+�/�ԁ{+�U�6�{��O&��4�W��{�ő&�CqzA��E��u���ٗJƬ�����s�>q�k�P��H���G��w�o�Y��]F�9#��� �5�����s�n��R������C��� �04�Q���H?��<#��sv�P:�kp �� ��f�=_A��m�T���z)dt@��ӜųhW�\h[6�6����)U-�j�9�۬��󗢇�r���p,|����`�̠q�T�,�`�?���*��n��di5fBR�W�> i�I�=�B��C�����ʭ����y�p��B�	� n�bg����!rE�* ;!��<�B�������H&��c6 �?�hrI��a^����:���O�c�d/�J��il����=���
�PŇ����_d�f�䅹;r���ND�?��NJ]*�ϸ���,����m �_ڰ��у�\�g�5��'����/�n~6?�pc{��O�R��{�nظ�jeJ9Sч�кcl�����:ަL�a��YS�8/�\Ĳ��W�lx@������9T`�4{�9�S�Ƈ�#�NTD�<gIB9��"r�T>���Z
V�5����OX�<��?i�|��>;t.��s���?^�`�U}�tTN�`~�<��S�.y%P��K�e�e�G�;�F�Y��l�-( 'Ǐ�P�UG�v�P���u�I��Q�J՚[&؞������C=�	Vb68�PO|u�p$�!$��5�\��Q矿���0�I�����""H�h��Eل����^��p�b=Ȁ;�q�z4ƿ����* I^O�����C3�zd�mӆl�����ސ�X�HDƊ嘍i�`7]h�<�C��*UK%3�h@��$�|��A�od�K(��ɏ�)�Q���N)5�y�B('Ih!h!j$�ǕM|�жi�Џ�7p?K�$��J<���3A�NXA�w��\� ��0�j$�}���$�37�k#̐�I��Åz�����G�\���7�-V/�[�O�l��'��{�%�S�&.�g͘�tV�p�����f�����t�+��ꡉ8��w��ͳ@-��I�l���<�8;�� 9N�{�����ϥy*�?��C �vklHY6�m�V/���ά��(
"� �X��Ŋ�3Ѷ\x���!L
�'I^|	�-�s�\�5��;���9O�����ij�e��+��R*{���	-G4}�ߛ0�&�:�O�2�/����{�i��D�T��o�+�����'/� ~P���N�B�#a!� J�@��G�'`K4�����B�CT$o�    IDAT=��5f8��'Z�����UK���֫Ikk?b?r��z�I�}p�͟;��1�	�EG�F���ybŊP'��@<8B�������AU/�+��{.��sm��טkY�RZ��ϵg��2���O=,r����CU�T�,ޒ-^0Ӗ-_d��P�Y2��`
��?�2��l����b��/& V ���_��C�dE��E�I�Q��a��b�!(T%����G
������������ng�O=���n���:���$/xp�RK�)�Q��G�"qy)|���(� Z@��(���Ђ밍�Y)"M�Q/�ŦË�
��[�Zo�I/�L�(�&V�ZKZS�D��/x�z�@%[�p�͟7+d�B�h�K8y\�<�-�08^�|@�':ģ�Ik
��B�P�gb=���2fEJ�Sʌ�tT���2��8Nk�Q�9���:���Z�2��%S+�<d���P���Lc�%S���<�*U��:�� �zb� /�y��Y⥈,�a���5�.U��AqW����x(9%"���g���K0傥����O�4����G+�P����h�l�F��S�jH���-t�pnii�E�e��,�;�vR�66��uF�5��Q�o�j�x�I]���v's��}m�����>K��?Md���d�}y�1�'��Λ�%��//�k8�G\����o
܉���\����X1��p4ro����}�=���ϊ��"�c~Jy��U3�O�����>��t�Ϥ�V*g��9f-�)�2�+18�A��ĩ�f�z���cA�S�z
0τ�=�aťpVi�Hi��E�D�Jm(d�L��ǒ��CkS��\�ԦN�l���>Ι��<�4�87	���{��4N�R���U���b��v���`��fO�m��_�9�f�E���MJ��kRH������?�I�#�H�����iq��+��n�,�pm�6Q��?b��<i�l�e�^�ө�QJ�'v�c]����gΜn��~�3F�	��|.�WQp�����_q�K9���@��p��B�3�����g����w�OQi���?3�s>���:E�-=��Z���� �C5Oj����9k�]z鋽�o2I&P�p���!ڇr�p�(e仼���p�3�T�q�?����G��	�$'f��6�lkl�0���X�ʢ{���?�'�[���B�D����Io9+9��K:WC&/N�J(�If���+^�r�0n�s}D��S�N��\2�0Ƕo��}l	o��%�dh�
� ~�EI�UGvM�̹t���JV�^��b%۽�!��M�Ȃ��|�7N�f�ut���&%~��U��G (!e$�׭e�~&?E�Q|%J��Z��
@8ʔU���� ��Q2���
�hR
�>�@�E���~r�X�6�(��CNa�<��!�\���F����I�o9�d��}�C�+�\t"�a���C��d9�"HX#Y����"K�<������h�g.f�]�|*��퓴B�7�wX�ܬ��n+W,��X-�h�bŒ���[(a!�����;`�&ݟu���6Dӕ�^���W؟�ٟ�Y�B�zq~ɘ�ҭjT)L�(��m��\��Ək�=��'�0c%8�����;�)���`��fa+4t����Z����ꎢX�3M~�_do|�묥�1X�>|�v<��u>hM�F�=w��w��:e�KUK�3��J-6
�!P�v=un���S%�M�g�?��O�#�xp�>��{��ah_�x�v�z�N�8`�B֒�%c���IKc�x۳��{߃6�������i>2����hN!*~�vv�u�ɆV�3�B��E	I@ոK��(� �����åB����G�5%PD��k1&e�J�]	/�[��響�
�IX*ƛ��B�{�:�k�\OUe��7����s�R��e)Ei���sܛ�Y��ҳ�7����SB����5�	�_O��~�O��P�t*f�B�mް��o\a�b�ҙ8ͳ<ο/�9�Z[�ٺ�<ڇ��yXl,P���Tۇ�Y{���k�[�盽�P�-@(P��o��"�٦t���Y�\�\��k����<��,��#X�����^!V�>�
�P�`}O�'M�r�Y�u�֛�{z�=S���$��y\�)S�7_�*����V-Yϩ���#?�'�|�Nv���f���/�bp�]�l��^��#` �������
�S_���ԽA�!���fΞ�%��4
�C� 7R�'����	�9u�N�<l�~zc�V�X�XC�kk;����Bm�~(��}��3X��Z�lF6;σp �pg�R߈�a�J�^�q�?'�U�+����Ł�����Ɛud>)��f�9c�GF��!sH����q]擒J����z|���N�Q�D �_�� �}d���&L|�^�ʳ�ٽ�AV�E�����B�j��{��� �oX�� sĵm|Iܟ�9撹C9�w�&*/j�L�2�+�j�x�$.�mP�_�Ϟ�<�G�����S�e�r[�a�U����$�����i6a���I�@��垓!䓤O/R*�y�k��G)�����y6�d��A������#�@Nb)3�I���K����{�b��{m����s�c�굶v�&���%�Le�;��fh���BEÿ��ugga��[?���s�3|��aH� ݛ�'o|�l����kk�i?{�^���MQ�b�jI�!�j��_�%KWٺ���9����}����)�P�p��+��~͵oqI ��<hm�G���zmr�U�=�޶ݎ>�!��$2�&ۻ�34sɖ�ݤ�ϬuW����q �ď?��mkmE����u��9�S8(<֍�u@�������=���T����>�`��6�8�i��e� ~��O:�p㾔� �ɑ@s�z����cԴᙼ�s<X`���Yփ}��!�(W�㟱"����������C�s;�^MI���O>Z!�{�Y�ʝ�	z=pO�hQJ��_��"�3.������X�p�wXc�\��&h �%�����5#y��O-�b��3|�}⵼��x�fM-m���6v�T��˚�.�֡�C2c���,}~9��\������;n�Az#�����9�;��B��#���<��`A�R�q�i{�ч��'wG�1�K���z�5���V*�l` g���?��Q3�a�
��{����m���~8�w����Z�Z�7��Ͱj�h�>���������`��KK���w>W���S��_��lŮz�[h �]9�2���� ��y�k�>��O;� ro��M�D�i�=(���?Z��Uc�I&,�(Y���־o��j%�P��\��G���)�?!��_�X-�FJ��� 	��j��@?�Y^��KD��h�<� g�	 ����e��?��?�k|��?�/�@�i:z���ŢMQ�N�� ��V��F��É��`.Y�@G.�=�3`]L�:Ʌ%�)����\��hX.T'eLX>T[���vN�̯��9�K�y���?�k����;4|@��`�ױ�G��P�Mj!!d�/h@ ����{D�QdA�r�
?t"�E��BbL������g�UF�}���)�`���Z��֭_j����9#0n��l����a�Q!��]h��D�F1���:0f�����Vk<eͭ-���WzIg�?���X��a�{�ö�\>�O2Q�#��m�欄<u�{C�|��kv���,�����~�-Xx�o��|ͅ>��|RZ�(�svk���?� �i��ٟ�ɻ��a��}��ٺ˭Z�Z[�.���]��Y���v����f�tۖ���9|�2aY�K_[�G( 	��}�{���ń�۶�,@��06�\ФG�},n�Z�j�y��v�X��k{�
���
�����q����M� -6�G4?ټ<�f6���ƾ�-Fh�@�2ln9����̛@t��j)@{�'?�@e�5Lj5�ȸ/��T��µ��i<���+!r��E�s��d��C��-娱�кyV��5�y��_�6���ͅ@���u~��<��'w� �U����b>���p=,�xz#�Rv���c��+Wz�4�{
���PE�!X<(X!������e/1G졨������ь��?���D�V.[`�6,��J/x�����Y�-o�V��{�s��sJ�y=�9m'=������s~ޒ�}��wT�,`����+�	�|��{��߶���)T�N���o,�Z��}V*Ǭ�x��ʥ/�K.y��3����ӳ�i�r���=��붭���a8��DC�9m��p���J��:q�~��o��e�������ug��R�ӝ����l����6w�b�r��g��jY|�EW�q�U���e 0���"� �5����DȌ�Ex&E���:����y�
�~�E��D������i�_����
�D�'��.~_��&��w�.PD���`i^�3���IVh�h����g�xa#<�3 >��(�CA3Ѷ��];��� ���}����چ��h� ����}$˫\)�8xa�߸?��3X*_�Hx�G�((��K_�VԞ��#�lX(T<廔�� ��Iz%�	j@����}�.όe�����)8�y߳k��=#�g>��\ ���G�T�'�Wq��zU�P�'I!�ꀭ]u��߰�҉�F#��Y���u�H4[�d0�Xܳ� tѢ�&g�g~���>Ŋ͘5ӕ��v�g�Q|��P|�s��_؋�S�'��c?�x�-_��&�c;v�E%�$䥬�7k��t���v�D����`���w{%�#�N:%�s{h�?^��?��������y��m7�`�I۷�q��[_����V.�Yǁ=�M�S����Z��C��ڎ��KVx�T �k�Q���w%�GQ��b��C�븃D����>�P�3 "pJV�����Nkk{Ҋ�^knL{)j�留�}Z_��`i��l��YV�~$�a�W\?T�ҥ��8>����^��Q�]8oh4_�X>80�<��&�"(&N��3�	���C� � f��C �e_s�N��v��2� &����ϐ�?��$3��j�O�<���������G�:S��b]� о�7_��^1����h�?/�A�#��cg~^��K��_��S��茙�&X!(<B Z뭩�ѝ��
A�傰Ta����������B�Y�*���N^T�ݸn�mش�j��OTi��V��9K��������4y5\b�CE�������hwkݣ},a�}�����7��)^�q,a�S�	5��X~"�9�(��{����a�2�8q����J�Q�L�-�-��]m^|��'g=}y����ߚ[�Y.[��|�c�Ѿo���9��O/�r�Gz�{�:��_�7
Y8���Ʒ��g���v�7���������|X�j%i}�y��+���w���e���Fʣ��������B��h� #��Vv����v���@�T��/9w��y��;rp���V��Rλ6���X�ہC��{�L�LC�
Xϛ7'���k����+�ꪩ�%����'������n�Mp�j<�g����;��w�P���] ���,%4o�V�Z"�`'�1 ,C�i�p�{�X�y��o��8��>%�X#iϬ-�`�<�Ȝ�7Y�'�{X>�=����>��<3���������+��F�0G(���w�� �N��Rr��ޔ^{I���B�OE�9R�آԠr:Ȣ B(�i�U	��8�D���c�#fӽ�?�\���(���O���[�fm�ʅ�y�*K'jV,����V($��a���0�����uʜתa�]!����٩>4�P2� ~ᅛ}MX�T�jemI�"�G�����??w�z�~t�7lŊ�6}�T{��G�Z�'/h���,�h��G���d�'n�L�����ܳg��&���ׯC���_����~�<�d��Fx������w��55��Z�ٿ��?�E�-m�W����!y���~��~�ʵ�=^��.�
�L6a]8�?��X�K.��M4/�M��p-]��7����nΣQ@���Wԑ�{T�|�������U�$%��*W�6n�4{��6��COZ_o1����m��6w������r�у��P̊� j��U恟�gW��*��h�\W	[��G��F���j��\ �\��o�D%W)�_��Z����
��}�[���9�џ�R�38e�)7@m�J@SG�~݋uT8��y�3��5ŕG�A֏��T)�?��b�?p�T��	�g!c�9�H$���O�mUP�/�BC׋�c��14���H,,�:y͝��N^�5���Ջm��%��o����:M�ן�1�&��~�R���{��J=�'a1����[�p�Z�I�я~�[�2.|?(������s*kN������g��g����1}�577Z{�^��(��T�1{�g;-�i��ǻmݺ�쥿��Ǝ�d�v����S�N�?���[g/��F�`�1aM��r�6[�v��,���ʀuu:���]����J7ہ���y脝8U�����\�����)�8����H���щ���ܻ��ݩ*f�/��hn�t���Ås�}�N�Q��s�
�>76���L|�����x؎�pb��Ϝ19�i�*pÃ?�*�#�s���f-j`E3�=Z�Rq *��<)��M���P�: #Z/��?@(�s}����=s����氢a�!�=�/�&��X
<#���+ˁ{�ys}�+��s�;�Sy�ų�󀇚�3V�����%$��3�¼���{pO�Y;w˴�V�,��ʭ���7��2��J�����ESro������i�E�:�Z�(���~	����?w�i��U<�w��́���W,؆u���-k���'E���%l�l���j�/Xn�\Ś[�?�Y�����[��Af���!jg�	��Z��BAOr�yvĬ7c���p��+���'-��B1�:�3ꊱ�-�c��?o?��Þ�՛�����S��w�|F����l@��Q�&O��K�����N�b�8�P<ekW���\s�UJ9+���c�#��Ȟ�ŇO��	ո�eK�(���.X������㧲K�����+�� �N��p��׹�@4�����pM����f6���-�g�'��b�ϓ�0)S�9�{o�=�}��lt��l���6s�3JZ�� ��p�0Y�d�8q�/���9p�lv�`����������9<�CB� �t��	��3C����4Y�(������*x2��a�������<BN<�����rc\|�5b�rƁPC�#�/������@ �(�7~|!̓'dM��kϸ���S��d�TB�H�W�>�a~� "�D@/��f�j�0�`��٫Ap�7et�������b��,C	,��>�KSԂ��W�N��ГV++Hc~
��4�o��L��^[�`�-[���P�������y���<j�B��O�����ʁ��k���k�Tj;g��r�-!(�=�S�e��Q��3�l��U�}�־�������',CK�B?��ez��6o���n�fkjn�����˭_�g��%dߟ�Uo�r����+>������8O�f�KUZj�<���T�����~��ֶw�e�h	w�,�`��۰��;���,.�@4HT{��%��F� ��c��M�1݋E�� ��!���>�i؃A5���=�i�|����!b�b�s�X���V,�(ڢ��'���5�>h�42�q��
-��w�r�g(0E���n����K4Q4~g���l�� a�1�e�XHD�`#�=959��4s��7�a0�����D�0��:"��y;D��	��B���p����0v7B�8k��e�#܈���K4 �{�
 �m���5'��H/�V���A� ��׮Q!5��8h��J��u�Þ�E�;�'_�T��@;���ח��U��5foHj�D���	0G�}$��\��=b    IDATG�ߟ1mz��{���������T�p���^��S�*�����z�2��6~�Tki�h�}Yo�B�x�O����H�T��Q�z��#��"�e@ԗ(4YF(6��Z�`Ǐ�����ܹ�:vX:�r��YҦO�iny�-Z��b�����/~�KFU"�Fz���?ra7B�b�@��@s������:�?g�d{h�`'O��G:�6q�T�>m���0�
� �qڢՉ{�@�9d ����w~�@�8��� p�1�f��gpͬ}�>{�G�����U�9�N��Œ�u"g���x��*U"�ʶh��={�����5���c�U��o��Vki��I���p��Y �Z᪀. �Q�A��{r��	r� ��L��;L�� �ѦBݓfP"bEEf1���y��Qr��/͔�� >�q�L|r-7���C# ̱$�=������N4"< |�|��)��%�M��~��pX�V���yf��1��x��rҨ����s�8\W&�0峚	)-eq�Q�_�蜨�XV��Y~}G�CV\0�0	Y.<{��s�����P��7�v<Q���36ab�ūeKg���L�<O�P*ٔi���/���4��>�XҊ����T"��n�5��jj����'c�p�����|D��(�2��o�iӧXKK�u�:aǎ���9y��Ek���lμ��L|���;v�W��ekko�Ʀ��p����+F,�������F�m��������
[�t���9-^E����꤀S��O#Z�*5ʉ���&�Xt�.g`А(���녺�.p y��H��fO>��>��V�D�f2�Gi"���\���{к{�Pn�g�3g�͙=}��	��4���Bp�]]�|��PG�k�dx�MJ�����? bM �p��������NT��ׅ���a�p1.���4l~b����.f6�:V �6��pFx`�Y�ϸ� �p����j��u$�@���s*�-���`a<<'�\�
Q_�����-%�ː=��QA8��9a��o9��KQ�;�ы�����×����t~2�*�w&�"�)?�׿�w��`���'F�[J���p ���,
�u�{3f̪w�:s=��\�ٚU�m�U�<x��$Z��^7a�]��_�^M�c��A��),2�����@_���;�|=�?�>�x�;˺D��x֐u�|�+��+�!(����l��M[[�z�Fj��FX�߼�۱�I����G�p���)��;+�}Fn悃,t��@�ĭ��j�9k�4��.��6n\ocƵ���d/c��'�w�s�k�Q�5�Iy��k��B:|0�OM��W��8sB=���u}��V��;~f'�z;G��	�DXa2����~���!��@ uP��ϡ�H�l^�3P&���}�k_qpE�E��	��xf��d0��M����{�s���3��X U ��2P$� n~"��_���9��\��.L�Do0� >Z5c"��sPX ��'z�g����7�@p���\!w�5�8�@�E�>'���Rh����>� �b`��;�[�M�	��H/�.�0@��v�sF�xi�cBԌ�'��Ⱥ�x�τP�rGi��>e,������ʘk���sO���@��B���I{e(D�?�$�,
B�4iJ��^�?�N��n��ev�5���Z*�L"c�r��u]�w6v��Z��� F!�Y:�`U��jN�p^?����A��NJFdh��V2�{��nͣ,){P��]�K�㖑Q��]I?X1w~�N;x�@(��sX��b���j�Z�2i�gea���8R�#����K�ZM��%�Ny	 b�d?y�7���{,]o����,8��& ���������h��f`S����7Ra7�:�&>}�����FS���������?��T�
�!�J:��q�9G+��a'�u��� �E��3*MV5  ��\xm �a�E����y�&��� ���=�@�= D�����YE�p-�V��=s��m�{@�0���	���,kD�Q2�@�]����@P��C �yc�h�(? !��"���hrMb��h�0i�\��M"�9�惤D%�y< s�P&"�u�>\ۭ�tz����9o��~/�c����S�eNX�B�����J��ҳ�I � Z�5�%��q�?�f.���[�������X������R5�i+T����-8υ���i�BD�"�����7�)��66X���^����U��^�0?��^��b��;��Y�g��:8�<�´������Dw��U�EK%C2�sWü��[�ʒ����C<�)�t}ʋ��J)$	ł��� ��kj�;:,J:�	p���x�l���z�'k�U�������$�z̳�?��R��d����;R� ��4s�8
�s�eL�P���b�n�*iH�N �h��zդgNWϼ�.�Xڧ�4F��84�����gĽ2~Ơh �3�7��6�h�pW��r�	+��9S�-�仌��Sa��}$�枊����O8a,H����9�F)���h?��C�� �&;���yQq!���^e}��e���~��{�}�s/|-�e�K��B`" �h7o?�:%X��	+,�#�	�G`�Z`/Θ>�����!bi(��鞵5+��u�\9Jz�k"��է��isl���ij���B�l�J���S�롞��>p��Y���&R)+�r�V�/��5V������"��(b�>7D#y�!�h�4��M��j}\X�����b�����}����
fR�%;���j{��zCo���A
>��,H����^r�Ձ֏���D��P�#��'�[>4OBBh�7O�<�����{n��y��r�R�c���p��u�k���g�?��q��(ِ��IA���<��m��1f7��|q�q�r^lz�I�աW��(��p99��:5�L9�&����j��:�-�V��Ys>/�Ut
ϫ{i��$%����D"m�46�����N}nDo(�����XO��G�W���}�;4Hi�DXae<���^��1 HZXS�?�+�Nܓy��}�53��דlV ����ʇ`]��_���,�:8ЙX}�M��O�0Ux(�+����^�2�X�X�Z(�i�C�W�����ﭽ��~���v�4ѨkV)V��e�-Y��2c=��.^iώ�z
����	sa���ߛ��S��\�W�d͘/�rg:���9��N���+8X ^&\��H4�Z�{^<h>�P���(�;��=�L�� u͟�^�����Hl0�������F�_�%^��A��g8DD�l��B��Y" ������ 	������w���Y��S�*a��G��͜5���B�؀����w� /LH�=���V4:>�Ӕ�D�h�p�p4H9���B��h)�(� 0��VH"��eP&h�P9�Q�T��{P2h�h�P��JEà���g���c� Uċ(\?��c��l8kq�)����$��1C��S���U/��% �B@�F�Eĥ�S_��9�/�{(�ZV�@_�������#掝�����_[*�v|��I��E/r��ń��9��<?Bp0��r(i��ի9�%��4�	Ʌ�S�5�2��$�h0�/�!�G�k!�
-���Â?�/��Y.{�6mZn7� _��&�*��]a��-�l�l���Rҙ��U"D�Q�Y�����ł��
)4n�+�����S�J~]��{�H[]���[ �
_E�Rb����>�����3k��^v?��CæB�?U�L:���o�����$V]�ߞ���۝�� &�qSۣ��{��1���y
��Ъ�{�d�VJ�`:�����'�!�\
�Ā>�ihy2>��������"�	�c���w�#4X��8�8`|0g 	�K2���g�Q:T�D��!L��Ǣ"j&Q7X]|W���h� �N�(�%�b�B���1_�7@d�h��;�	�?�G\�U�q){��8]��'m�>J$����hd�?���_�h�]����O*�27�?J/�$��o��{q��g�x�R��pt{�{�A��G2�`f.��TL?���Ǉ�~�~.��%N^Ԣ�!/���b.�k(I���6uZ��sZ�W�o��C���/jum��/���J�d�r���/�CQ�������k�p����`�>)/�m��� {�hG�Z(��K�'�Gđ�9$1h�`�����?�_q����t��ax�B�Y��/
8/S�τ$�@w�0(��
�BY4`�)�C�Aw��������А��0�5F���@"̀��y܎�g�r�A�fko��K��J:W-4s��l4�_�9��V}�e��1���o�fO�����I�*��.��E2�J@��U�	`��4����@  ���P�8 �d Ѐ�*��|�*Aa5����c�!��.�
����3s-��  
�@�po��8H8�X/�<'U������/�3�����%? �$�ƺ#���!�g]�2UrӾ������lf�q
������Z.�����!�%��ĺ!�A+A%`�ܱ�]�/���|=��L����^w�y�3��ZN��
�cF0c�!DP0X;	��t����N���ok�.q�'Uݮ*��
��ҍ�_�zMj�s���רµ�C�p�cu��c%Z(�U��:�pܑ�߱�V��7f	�r��C�Qh(Q�N&�5pf�0Bԋ�&O��t�nݶ���==�?#�ӭǝ�1��s���>8xc!
Ӌ`�D�������%�@��()�;� ��h<����9|)���1^���v��n;y�Ò�rp�Vj�H5Y[�Q�羇O�%��?}����f�h�`0�n�r�cf^���ޅ  �s -<?`Kr?q ��7MH�͠�-��`B� ����E�>?4��5 }�w��� �.s!�8�l���z�j   �3r����h�|������R ��x&ƅ3ap	 �e H?����H��b P�)!�b2>r>��u����c8w����A���Љ��n!q}�A�s(�J��Y��,XM>������M����S�3{��W��khl�<ւ����{���G�����SXŬ#g��V��8�6p'�+��Wm�t"n�j�V�Z�߄�-��Y�Hᴄ5��n���Vs���Eע`����{0;��\{�gF���r�d[�l�$?��9�Bs�$�%�	qbSB���P\���$!�⊻-K��fT�h$M߳�>���=�myfd$�����5�=_���y�zֳ���փ���V�T�-TCX���gT�O��H �;FX���k��]r�O-�/"6 ���Q=����ܲ��==ݿ=2�G:��+�y�j���@�x$��[�lSo��2�'+�>�>��8m�U���ΟI0j�7V�C�vX{�~��=f��R*V),�Գ���n���������o�h1��gW��@ �D���-�' �{>t���j�i&�B��` �X�o�� ���%`�#��^2� �=��my6� ��� e (�}��z��K�P  ǳ�;W ���� ذL�2ѯciC}@��?1�U�eL� 	m�c�i�6�jG*.Yi���:�����^oL�PY�˟g�j�Pb��.�ω�	�b��b���al�� zyg,*�w������챋6m�׿�j_t�&j4�+��Ip�X�;�U�s��Ρ5��zO�w�����b�}y�x]��9��G4��iy��3��ʝ�Z֊�-\��.^�ROh�z�c�< ��w�>��	1�x�p`~�+��@��lO W�cx�����%@����޳����0'��6}�uw�z��O����G]S����+7o�FOo�F,d^��C���A��� �Z�c!1f�R�Z&I��t�^�SBQJ}���A"��5X ,e�q�'�`��g���^��XC�E*��G�7��]?��r��54R
~v��uf�
`F��k��ď>��SX� )�\�pŽ1��$��X�����R�@W���X�⻙����o �����Yx�G�`����c����B8�TAE<--tx,&PB����|���|��=��k��N:�X�B'�����bժt�(=��(2�O~	%��p�\�!��}��]�Prܧ,�����m�\ v����x2�#o��1�Yp��x�|�G��:V1��vIlǥ����546:��x���L��њc��1�v�{��Xg�#��! E�ܹ�O��}��O)f#��_�ފ�~�t:k�r��_J6n�$��%�Y�P���x���\�Q��$fG�/������|�j�:v�0j&�l�H��w��H-;�~Ľ��/`M�'#�y�hL����4�O	V����O`T�g��C�\(\�B!��{�sN�v�MwW,M�5��bV.Pf��_���f�^>/+¥m(��J�*H'~�c`�B[ <E/&wb�v�c((D��'�T��6s��`����G���~�|�q�>Fk"\I�y�Y���>:�x�G��������P��{Խ���s�9@u�X�܋��`�K������<;�����m$���`���^������ه�� &��]��K����]`aSo ��V����X�ܧ�`5����R}�����|�uJɽH�X|����"��y<�2�B��NUD��2:(+!�G&�;�
���/�Z���b��Y�y�P~|�u ̞��N�9�'xx%ހ��g�������ؑa͢������~g�w�9��g�s^΅7�K�ϙ�	�ּr�	ڧųy-V���,��kVZ"R�����K����[��l��(�� ��k�A2�����Ywoh�ٟ�YC*���?�Y����ƻ�~��+X�q��T�b����p9���?��;��1���>�Bry���UJ�S����ӯ���ۿq�Y���>f>��������I��Ix����CB
3�$��E��
�(Z�e�B���=�����h�W���p�'Mg�Jɚ���)cbx�-���v��[gW�����q�6f͜�Kny����Ț�Z�p]!X���y2���r?�G� �~��@�y"���z��"��ZM�	�D$�H�TJ4��$��p�s��¦������R�<�)�NV>����<₹GY{R�pn%�q/Ҷ�K��O%��̉�p���xMx)xP��TO���[��?��g��X��t�L�����c��b}:��#q�Jc�w}��>|/�������,�Jy5U�Z����� ����dB�(�J�8xW���+?���*��s�8~����=�W���6yJ��k�>��@\�x}���{m _�δP�d�¼L�k#�u����.������7_�ޗޫ�5׍���Ҽ����Պ��q��/���C"#�9*5�ϱ25�*~̐�w"?`���c��vr1eAk�c��p��sw=�t2�I�:���e"���y���
*k���$9�8MMf�����V���aY���:X̎v���V+��Y�Z�bs��O0y܄�6P(Z#�,zXT��/�ksg��C��h��`�t�LƯ�������
P��1 ���Ƶ�>���'H�*�zЕ�㗼)q٢K4Yd-�2Q� xn���6r���i��z�N�,�kl�V�����{l+jMV��1����_sl�A��������D�������Ρ�J\ �
�'����*��#N�	����,f���pn-bl/���#!�/�E�k�Vc;t�X��˟�2�C�"���7׌5;�F<K��<*�w$�oȦ-_豄ap�,����2����%2Y�4�;����N�����U+�iCRk��ݻ���@��\�x�I    IDATt�E��>��Ϻ�#��K��]=�%.�-�m��ܠQ�o���E_�~P���m�q0���ij�X$�6�yG�Dj�k�{�m�Y���}"0�e�9h��e˫��=�iC�,/�� ����yйm�|� ���-�1x .Y��r�ha�� ���@�i�X����n--��ˤ=��#.Q��g�Z����{i2�I�d���ϛm"Ji$��m���+� ��T)�p<Y��U!�wՕ��U�&�����_]� �_�qh����\T���������-eYr�L��D5Z��S�|��k�z�K+s/J���U���[�eK֠�x- <S��v�8�<C DupD;r-��� d@��>X������N��I8�Ȇ�������u�ߺ�)���ϖ�П���w�x�AV���<h3f�t�b-��L-Z\;�t�p��"������}�!�����G�8O�:#J��,��v�U=�.�i+V,0�-���܍��GgL�n���ם�)�B��x���/�r���h����-�_�ީ�o��g�3�����_≃��/hl8��lC:�S��J��?z����$>��9�*������?�Ο`�T�o �믻��]�B��\���bu�o�ץvP��;d�q�A�z��]�jչN��8TO�>��q��yˮY��Cf�iY�X������c�w?�%����)ƶ��_J.D�aGfB*8�X�ҭ;���{����e�>D��,]�O&e-^�ʗ�{�uC UqY�ҀkR`�����5�-��N �`. �w�EO�k$�C�9��L.��J�d�s<b$��4��c��*�>x����y(%���Ȋ��X����5h�g�q�d�s\���E��hav�2R��χ*��Q򉡼�
��=���r���=���s�<�V�ȸN&��HB��3����1u�+��s���i�?�i�S�Ѕ��r��p�5�x.	���)�0<��S�k���Vڅ�s��{�� �$V�Ž�������K�a�W�������@<�"���&��1�������[�t�0����cbC����pA����d���t���93��<���E�u�ڈqv׏dw��c���b2u�4��?��$y�V�b���NϘ6�9t&���|�2���O����x89
�o-Ł���y�L�@��Ǫ"�&:���@B��A���B�`;w�ԺzY�B����>�����ms���^�9�o�J��}O��W,d��:�Fp�[Z��D:��2�wJ2 �h�YXP��FÄF�$���Ft饗xP���}��>� n0�8X$ @*Or,�E�)E���J�.��a2�h��"�Ċ�o�&19�2��*��;�����-�<=p������Ce�M��Y9/|0E�xތ��	 �x�я�t5Ǉ.Q|����F &c�w�@8cL���`�h��x�=��� �\Ƕ���R�s�����B��9��do ˟�� 7Ή��kg_��k"������c�?��յ"ϲ~���=�l�?b�;рıh�T_ۇX��z�{m��e��5���v�o��J5n�R�Ə�l6n�r%�u~��{�0�w�g`���_��7���j�f�t�����"��2��x�4|g?1��1����@��qD:s���y��<[�>�e2$�%����=_��sx�!X>f��N���@�	N�>���o��V�<�]�|�߶m�x�>;���z��2$-�M�.����3s�"SU|6���4�L8L\H2 ���f�Q�< �Ԯ^�[��b�wv�ֶ�V��F�5_�5��%�wo�=��v��F��h���7o�!۱�h��y���C\�	�\'���@� 90�lQ��< ���H��&�{��# �dâ�\,,,"�+��)��YЋcb9�|Ѣ�3�X�XX)�`Cͱ� �(^H b�}�+Ã�<o
�2Ӹ~����ɽ��&.��<�7����ޟ㑸�+ә�)S ೨�����=� �����G��F���2�E3��L���ճc�O��O�y>��V ���?���?���YE�?��sƻ�9S��g�"I5 �3�(����wd� ���q����T<ԓ��k���˸`Fyĵ����YWح�����X�V����;$�H�$%�B�����l��ɶp�
Kgm0_v#�󧼇u���4��9d/O�1������w�B�\�2.	N���sc�+��{���x�믶���pgg{�=�����S[���7j����k���um��3�Z�y�����{DQ����=}u�[F��|�)�b�6n<�^�ZR�y�kn�k=|���U����)���Ҩ;oG���ŗ\��\}���I��Z�b�P���L�s�� �﬉	0a%���j�hR��ԋU,?pܞ����
��Ɇ�Ka��UϿb�X�-�P��U�f�(�P��)H��|Os��

���ʱԙ�ߋ�@����ŁkYu�yVX�,�,xz������aq� K��,(���� ��U�p�u�Pٖ�3�Ylx)�6,8�EZ��]�=ۯ
	���\�!����,"\ 1�����0tV4�b��d	�+d�+נ��|�'��C]���b
Xq� sWO�{9�a�0f9.ϗ�Xt� �� c��v|xWlG�>j�o�y�8�Œ�(�8k.Ԃ%p�ߙW�'ȳH�����1�����_��������v�R۰�����K��l��6}�|�0~���|C�8/��s�_԰�+���}��N����*6y��B�x~����R���7�)��*��n��6��?j��6n|���Z��>5{�寰Y3�z����vo'�{S<��8�7����nX�����k^s���a�%beoܞ�Ĭ����=�2J�R
���{��y��b®������L,'��QCrԣ�k_�]@-�D �Ky��'�?n�Z��F&`��e��n���\*����=d�����w0wsm���,(�H��������d�2��` hi���bun�`u�`�tx�,�,?��9�� �����>@V�,,HJG�i`U1��o��(րE�D0��(�@k��%p?瞻�3}ѕ�;�Z���k`q���Y�w}V�g�ǀ��҅��?���y�O�p�Tw�= ��
� �Kޢ���G��R*	L�N�g$�'�<��}d]C�K��s���ȣ�X�޹>���'�%ZJq����}�x(|`����y�#.�{Q@�,�������3�k#�>��_���y���J��n՘M�:�V�y�������c晐��F!�9i�|Ǽ��_}��LG��l�Θ�)p/�:�Zq<��^���&����֪��m�Σ���v�Z;�d���Eڑ�.+C2��|�M�8�b�?����n��.=WŉN��>�7s!����N9���=�o�tܲ��v��mͪ������u;ׇ
������:�TN���.���_�T8@�)`	������2�\l,?TG�v�$��W� �Wy��
�Ճ�J�j�׬��նm}�ʕ�gf���}�?��J����"/��?�#����\3Vu6��4�@������p\,y����m��� :�29��������"l <�?�����e�1�U�sJX� @̢�����n�kp��_q����{-N�3�[���11���\/ �W�g�f%� �b��xlâ(�7V?�f��9.�ͳe��&2��3U��.�lx7�[ �Y����<S��8d9��c9��J��$�,2�I-��s�/�c�O%τg�"ʹ�r@�f�xx�.��=��5��X$��)��:��Q���@
,�ݜ����;Pw���\�qKe�֬Yj/8�b������N�l���h�:+�Vȗ���?���{Tq4zG�I�P�ǎw�_�t��� �����^�;�`Jf��k�^�f�C��'�s��J���wYC֬�1c��^�� �:�I۵��i;x�î��[v��K,�����[n��C��zE`=tZ����C��>Κ1����m�R�;c����.�� Q�:��A����~;x��
Ť=^��3�z�D& /k_*^
r9^:�@%K +x��+\Ѡ@�`�:`r�^Փ��[��X��a{wo�d*XU�.����'�)���ޖrΜ�/��~��w�&^�g���w�4LN�^Ԅ�f�� � 7 �}�Sn�����-]�@��W2S�K9�&�hY�R�̤��z?��z�����-����{��e��j{ (1N��Иj��9�ԓ�e;%[j�^χ�=�
���?��8���zO����;������ ���H;B����kd_�)T(q � �Y�J��}���x��w�޾�6]|��Gx'�>X<�b�|����g5����jW4u;�x{Jv`1�	P&��P���%s��;)�����Jm�V�^b�?�;y�����'m���6k�Y�m�b�A�Ū'|�H���Z����j�x�c7�ڇ�>u�L����s��0�0Jx&�R��ϒD�K:l����lŊy6u�$�����BE�*I�q����=��6�i�����u����.>p�e��[ Nk�߼e�{z�Ӏ�1d=ׂ�ꬕ+�k�bM�������wϝ�i]�r�==]��SM�u��:b�r�����.r��������I�t�r*2��v�%�A��h��i"^�R��v�x̺��z	
� Z����t6z�Vk�h�"�3w�s��:��_)� ���I�A�,T~�"����lϳ�X!�: ��.e@*�\���\+�	@5����� �&%?9�~��nط~A�5�'p�3Wb��Zt�VO���X�ܯ��h��4.��K�(J�d�k�X
 �3���g�������pmx-����XR���Y�Q9�!��>ʑP�-4���1c��9'@�5J��R@����� 8cZ���?~�����&��H��Ϙ,
����h���N^��_��=p�,��VZ2�j_�z<&N�yα	�g: �C.	��D��D�% �?�2	�֗��dhlø#���Ž��c�|b���!����c�����b^��ҙ��ݷ��w�_*F�J���iu�����U��� %�@�홝;�ٌd�������_���~$�'��@]�t���~�*�A��;f���U���-�(��C�^��C��y���Z�Z���g����6zEJ&�� "V�^:?���I�$���䤙|���0A�(�������jǏ���������K��V�V2�4��t$�t�Yͻ�-��_��{*��k�v�zB�Aq���J��W� ��7�&)��ǩ�(IJܴ&���kW�W�e(p�'V1ϟg+�M��.���7ā�� �R�7�=��^ �u ���s~�'���iw}����u���&�/%�AaQ�=q��C��/���
���g�;��' U�`�B�Op�hX\�<���Pw,4,.3����q-HCG��Y���P2caN��;���KGa{��?���\7�� ��{�_�����i��Ӟ�5`��.�u�V���Z0�bi7q�e'Z63��.\l�Dƻy�H��:�hL��;��En��a����~���Q��������;O�4����-����]v׿��F&����{�b��Z�P���n���$;�v��{�?�J$�r@/�ݿo��3#����~�-'��t��9:�G2���'؟��y-�L&fw��5[��L����4�Vн�VM[_o�Z[�Y_�:��v���}5g��+c!��y�v���p�X����#L�%˖�%Ǥ����'���k��y�+���[��m��K�,c��7j�qaSm��N���G��)� �Zd���hI^Rp=^_<�:�Q�A�l .�τUr��tU?���J}kC�� 3�����A0y�K �v��n���@&zH�E.�ߎ��f{BD��[y&m�L���ST	���y�,�sX d��3����8�8}QW�^-,</>���#cDIO�PP�= ��P=�G�t�{#hK��uk�V�<<��<c/}��\����ze��3�ga�������o�UW��v ��?ng�\��@_�_������PG���3�S�$ׅ���_F�F����?j�dS1/�p����a��V)S�'��3$<��Kem\�D�p�ž ���&"����X�c4��'<N��/�ߺ��.@`� �g<d�~%��%:`�C�}�uw���i�N��q	g�}��/=a[��D�юu�lٲ���o|�Wm?��ϲ�H�s�� <�
�}N[��rOo�5#Y���2Y������k�s���-�(Y>�c�����e���LZ{�1k9�a���]�~�Ox&�*�r� �,� V��) ų���z�5��f"�J�+`�`%ԫ}F��#͖��,�1��u��ke�;����;N��e��/=|�J��fd�g��A�@8��]���� `���}q,I�ا�W��z�XT�J7��?E��L$a���(��}�p���H��[uQ�e-(|�8�hyql�~,`��⟵���!�h��`�����t�1��la�S��\��L��3Bm�3c�I1r�w<L�	),V+�`qs�LxD��.q�ߑ�@����}<+%)�W"�}��@��(����9�#��|���'�u�E��	�s�:?Q\1WD�`(��G�?���p��IXn��6n<�.8��}.�z&�]��U�)ˤ�s�Eό�{�^껇�����n�����qp�����]>G%&��ȳ��"�Q���=r��j%o�>m���HV����/b�4%-kv�h�5h��#���׽��]�֟ŝw��^�H�^������vǭw|����O��F������s�J{ӛ�h�j�*ł5��}{wz5O:��=�#��r�j=}�6}�"������PP�0�Eo����pR��A��2q�wדg��T\B$�N�T����	���
Sg春�p�Tm+�O&	�M�&[��#�u�;ޝ�Z?��f۲���*.$����җ�4��s/Ǿ��<���Tő��JR\���x,I,�ƢW�5��Q������U�< �X�Pyj�V��%/�-���5�/����i.spc,�47��.�l�_5� @Q5���m��F=D�`�J�����򈤢��&�a�g������έ��/����L��e��\���[s�7;�Y:��{��)��Z>_��	�-��X��={f�{�Y����<��cV�e0���e/}�{4ܣbP,N�w�������� 7�Z)X��xd�7EJ��
0x�i��K���k�T�]v�+���,���v�w=&�4~¨/�����?r'/+�X(���dMM��7�ٖ-[�u�a\�~j�g�>x��ʅA�t�B[�f�-;k�uu��D�7+�8I��ݨ�8���bB�
���:�k��+�í�:��y+7e���C��eqf�@Y@��i���5�B�xͥq����Ŋ:�c����_�Q Ɓ�J�~�,}��Jn+M��U}(Qr�)�p����+�l o��@ � B����j��n��nbN@�a�@7�v�;�AX�쫚F�2�M&�
}���L�;�ʊ����y*���o4�w�'��b1gMM	ה�� �{2���Ǜ9e�91h�Z�-j�`�s���Q��8S��jN�U����_��1<}�J��ŋ�Y�R���G�g�v��<J�'����Xn��]`��&o���Νv�Wi�EU��˿蜧5�o޲��{z^?���A���6A�3��3,��Oˁ����a�r��Qyoά�6k�\+US�8n�[Gdh�ؖ�@���ѷ�V  9'.9|,�����p��s�d+�7���ܼ���v��ak���L�EI�1c��+�c�e]�F!������ٳ�����\�,�_h���A���׌Sh@�PG0� l� �
Œ�Øb�3�P����L�|���Ǌ���)!��Ʊ��}�    IDATd��3( ��İ��U<�le<���ù�sa��	��"�˜!&�, �$u�D�wά���'(�V��8�}K&ʖL�l07�q�b��U�����d�r��ͯ�T��K(P��A8j��"������e����K�͛�h.�u���dA�3���빱p2�7����	�m��&��hs�Tow���y��p�*X �v�-c���_[{�W
�Li�<�Nk�r˕�����G��w�R��8m���nx�M�2q��T:�rp��8�b�W�����\+_�=q���FH~�}�IU>���KC�OQ����/�=��ּo��ckjL�@H)GFa�={ۮ����������,���&U����_�q�}d�364���+ �$hȮ`3c��R9 '���n�ɍ�N5�H������C����!@����>�+�CX��`�X�ϖ)ٹc���5�qCG�m)���I1?�@)fS�aQ]R�)����Ϝc�z����n��B�l���v��K�j�ު�bE =��gΘo���׽�s,Ny��d= �M�
�>G�����R�7_�V{٥���"o�k�:QAAeW�9�]_�}Ӧ��W��M�8ޚ��=������;�=��*�g���]{��-u���V��
ӧN{�i��9�埈k�I�Ʉ���7a�xzQ ŭ��D1Şsv׏�vK�~�,�X����[IxA�̠Ɗ���2�ؼp�1b��8J=�������ÛTSԍ��Ɔ�[X(V����~�����4�F�������w�������w4�7�lKD��ĪG#KRk�)����θ����PQ&v>jdþ,���>�O���� ���9�Z��k�W�q��^T�T�q��it�*����?�w�aI��
A�#`��QI�[�ϭ�Op7?�kk�[a�6��Ze�j�UJ9$<V��l��i�f���ן��x<.J>S��8�;��٧����3����߱��\ڍ����9F!:h6���ޕ��w������gKsY�	�%�Ugj�������:ފ2�k:ʍ��QhdS"�ͩ��
Or���x�R_�\�[xJ�����U���^�X�r5>�w��f����/�8~�%Q��!����~ ������]��Ԑ�d����Z�&O�a�w�;|���2^�%Ȃ��NYc���Ͽܽђ>@A� �C)�\X��we3��A��Po��Fߗ��#� f�U�o�Cy�Mݤ'�x������Ko�tz�H����]��M�<GEtǠ�%	I��E��C�t�2�z{{���O�
�# [Dȣ1�؎E�Le��� z5s)נG�����e�ןe]x��}������U�I+�)�7��n��-��>b��������K6��9-����ɖ-Y�^W�ҌA�*����爸$��y���z����&M��m���m���~�۾��t����à���{�0u���{�m_;y��:�o����a$ڇ��In�/���χ��^ld��ł�=n|hP�T��g���g�a�A��EF�/^8ٗL&0A3,;t�X|(%+�a8�?�붣GZWW��u
�T������.����>cV,T��3�r��NA�i��>�\�G���� ��3�c��&"��J�%H�$ aٓ�Ż���[(E�( zz����F���L#C���F���#m���,]�؟8���N����u���f��Xx�7d�/@!�9�^��zw�(ܛ��p���}�h�o���]�ܥ�I�?m˥�%��mʴ�6q�6u�l�x�Ű��U$�<W��p���_�B腲m�t�]w�[\�D�B�c��k����T]&)��d�޸=HxQ��B��,޾�^����8NC6����YG����X�V�O�>��;n���s>�=��ӨŇ�������+��O |�{h���Ui��cM�	�y�*�'����PJo{��<Y�	"����8zsg���K.۳w�l�ci��5ҵ+f�-�v���@�!��4v\R��5*�h�_,<�r��{V� �]C4���
P5R�0�@�` ���ᝳ?��{d�����V6��ˌ���Q�A�@]Я�r~���&su���A���m����!����9�z�=�}Y����#*U�^ݓ��|�袋�f.Á���s�]bm\�%�)�H�V:3�.>צ͜�u�JU�� �Hy"�'yEy,T�$�듟��Z���0���?�C�Kt��xv�R�@��˳�=`4��;������a1�ܳʐC�])�ĩa2\v�� ����Sq�/h�8��Fo�`�EE�"-���x�dM2y���O�#� ��=Ǻ��Ο	�d���YC*i�b�R�=vؚ�m��`�/T��7�������T,A�o-�nՓ�<��>�k��Ac�?i#�O�7��L����"D% �ÄfxY t�P<:�<	�m۷{�0�' ��l��>ۏ�}��ӄĵ��2����#���k�������V�^�F���G�g�>x&j��v2���`�?��J����͘�6��[��x�b���[��9w��SU/���x�Y�h�Z˗0�2f���d
'���)�h�nN�,��������k|��dqkjhp��8��uq�м,�F.�� 	��àO,h��GH<�>p�ӦO�����O���WC��?XQ-���>'�?�(E��cM��S�f@��M�H&��Vw&21QV0iFj�k)�,�IXS6fmͶw�V���9H`iii����r���' �MM������g�M�集
�R�@���ˇ�i�9��rI�b%3��� Q5O7�zD��*�xa�3V��?��%xw�I ��A�'��A��5r}���#g?U����b"��}@k@y��T
פ�o5�q��lq��^؍���f�zB���yk����˽��}@ۅ�δ�γB9$m�jP>)W�d���[�fNd}ui�O}�Ӯ�w=?%�*�ސ���l�G��u�<���,D;ɲ�1�^�e�{{z^7��_�h�jH��S��:�w���y�b��X`\`�9$e�äQ���n=�:&�Aޚ��{��J���"���J:?d���	�f.�梪 �<F���������󢪍� &F����82��� b��f���j�˂�*�e�Ŋ�q��1�����R�c��/-���5��kb��9�x
[�|�&F%�|��O�Խ����	>��I�+���E^F
s��(~W�!�9s��U�<�Ua�lM�[�֮4��:�SΘm˖o�L���-Rޝ���ۆ���%T,��{�ֶC�ٿ�,��bL<�P�d���r�(F#�&>G��O�8�� j!;�9Nw��;==��}a�����q��G-�ݯ�h�l3a�S���	,��ކ��U��D�z{�[_�u��Xww��#��-��v/�ݢf.���cD��⎁����5۠�/���2���]��ϻ5�A�hJy���Ϙ�8.��sw^���<	�r\��0�j����� {�(�r-c[Mdؗ�p�x'�cK�/V=�\��U�f?ߑ�����:ߋ#�~� �[��o�?��:Q��|�]x�9v���Z����x����>c�M�6߲��4N�B������s*����v��_}�
Q������K�+�K�bj�=*3S/�74���TOp��_��� �#�8,	ύ��~�Gp�Qd�);W�
c�KcA�Ť�����H=�X�i���f/�L[8�QjU�L������9m���#�왡�`T�v����?a�_=�cq׃?�E@I!ۡ��~�; %�q�ō���
Ń��lT�)���u�b1��(v���B�*�5J^T/�"�����!�W�R�;*�W)��Iu�D ��y~G�I��\�ߓ���������S6��a�
۰�\�T,���Ӻ�h�����V�m�}��P%���뱱Z�z�����?�s/��s�e$*�������Y��Kp��8��:y[���~M<�8#��u��~�7��O�	����?/��	�	��9y��M�ădo��*����:�8dmx�#}be��4:�V+)��l2d����0�Z��]���W�VP��?�\/]�����ON]�z�5M=�C숚0d�:hᡂX�
�dT�w��'?�I��_UQ�i�"�KZJ-@��2b|J�L�d�q��|Ϣ��,>��1�@U�gScP��XD���Ăǵ��S�d��x�������[����U+��mݚ��s��a"Q��W�	/�R��m℩v�K^扑P?(�<W���Я�q���J*��� ����<s� )|FYw=#�-C���Q^G0>��"8�;n����Qi��_��
�ؓ���xl����Rɪ�U ��B�8��� `��j��J�L��R��j%�V󖌺a�g2m�f�����l�R1���^�(8c���	�����>�B��,jh�C��G=�g\�DH��Ģ3�yM�9s�G?��� ��t��\��e؇r�xxT�e�����g�{�g(���8 ���F�-�	E�ꇅd0�?$v�����im����4�q��\gϜ�
�� �TUO���&V��m͹Km��gӧ�ɚ�g0���\��,Y��ZjF 8����[���|�;߶� �er����Ӟ�v�~G�GGY'�.�8��<�>����0����N�~�wo���O�濽���|�K�Ї(�@������Z[�ڑ�W���;��L��R�y�ZD���D3Ed�{�1 ?g�֘IX�4�HH�'R���ޢ=��6�Xƕ�R�-Yl�����Β�����&�#g�� /T6/�.�'W.�A�( ��Ή:��/2QJ%3�<}j�6���>�5��h��泟�ĳ�	�B���'@�<�*����8@�)>`�J��liJ?s�|��͟��,Z�9ǎ���-Y��ҍ��:	�C� ��c�P�͚��s��k ��j�����p�;k��P�V��,�t.��۝v�����~D��'��'���=P���l��[-z��x��>�/��)��܋�BA�u��[&��� �L����+7o�VOo���|�V��54f,ח�j�&��uM'3�
��i��fuB�����ِXLLJE��sTkE��+�<U*T��x�6����'��9f���V)�)`Ԝ�,W�)�,NF �A-n�.��s�vq�S|���:$9Tp���r�)J�׬d�_Mh�տ* F�H� �s��l���7Nd)��T^	�C�|�!���`��}��c�(���7��M�|�9�dYTH.���Ch�hu�W��NU攬��J��C�������?�����"+�������k�xUO,�Pճ��[�f?@���V)3��r������M�5T��S�[n��ٌ?��ɤ�ko�굽h����\�/u��� ���}�S���� ��5G<_.xŀr��� �΢LǼ��;�rȪU����`(I�ChH3�紶�GO�%��j^��R �d<e�]�R�;g͚��D�]R���b����� <���pl���冻����RkA&�5���C=�t"�T��;����l�\o�%1KE�Y��L���~���4�f�'l޼C5R�����I^����=�3������>��Ɉ�x�_}��սB%�i��JU�D*�ႊ/Z�e��y�O<���a�w��.6 Q�3���M�8��А�_)�d�B}�������F�-�xy�{�;$��PB� ��Y.�Г�8�k�
�˸Vj�qȠ`,O�:���s��	���P#��ڄ	Y;c�xKF�J�B��b%���[`/{��f�z�X
��q&�F����t� ���T&��	�x0ڔנX�EmK�Y�P�!es�Rq�l;�앎3fd�!���7`;w����l6m�R��r}��~#Nk�r˖Q���p��usή����y����'O����ϼ�C�����(����i���z�������D��FI^���5�k$��'|�l{vo��{�ZB�M9����T�|f�>{��m��M㖬��;g�-Z�0���b$����M�uY�xp��p�yNyB��ū�>/�	8������s��P�����ࣨDIe���ܵ���n鲅������;�UvA9c�����[�h$,S�%X�x��G>2T �kW�k;�:�Cc�{Q�,�(��w��]�HhA#>k�[�p~���퓌�N^_Tm��œ%[y�"[�z�{�rɒ� �4aǘ�4i�m��+㖈g��o2jd�blE��찏�|�{|�����k��z1�H
ʜ��G4\}�r	.��R���mΜ�^��Z-{��kjj
yh>X`����8�U(���T9*�=� ;����ͷ�t��i$�-jw'�Y*�����W��[:2�r��^%�h�;����O%A�ep�t�'�����A4iy�������+eȜ�J�����^�:.���������'��6�f� )��2��Fk9p���!���[&KY�͝7�� �.X5�s����������n�C�!X��5�d��A^4��;�6���+�:E����=`-�d���J��������c���a�(XI�h��D�W�,U;�Ia�����իz?�C�� �9�K,W΁�c:�V�7d�3�Pq>-Ķ��\%OX�Tϟ�>sf���z��r��֯[i]�֬�w�'�(�X� 64N��7\��o��P�Y�3��vx��ԧl0?���^L���8�X�'`�G4�(-l��+^��v�K/�d�R,dq����~2�T��=r=�rr���1=��\!gY�Y��?�W]��+��=o1�KE��)o�r��+�寸�z��z��c�;���O?��4M���sV���o�q&{���R��LQ;��XT
�s�Ԁ?�1Oaokuݶt�X������;P��С�ֲ�U���(nc�ۻ�m��O*M ��<���#p	�U���e�SٝJ�g0�z+d�X$FRA��x�3�:�S@ �PGG��h�W�,��� ��w��k��G=�K��:(�DUZ�	�sϪxn��f� :�?��O|���:������+�Я���b�@f���y�{���.��8 j%Ā?qU�9�S���D'�@�b��X�{�!����q[��L۸q�����W=�Z�ĬTIZ���I����.�rm?}|�ޛt�-�,�RZ�����+(m����K/���Z���ډͰp1Wd$�w��K.��z�o���J���ჶ{�km=d{����x�2[�t�-X�ĦN�IPK�����py���S���:�����v$�'��I��5kV�u׾��zl\cʛ��w��F�L��'��JO�\�
%���앶x�
�\H�ԜEY�L`$Ȑ���CC�[n�ś8��-o�^��eM`�SO��H�hW��9ܺϊ�ǭ����./�J5���mv���Ya��/���m��%6�l�Jb	��4�*p�:!����� rq喳���LX���G������f<�A�99�+��h
�!��{��?�f{G�, 	��$� x�y��\�V����Զ'}�R���BQ3$�\=��0d��/@H	
��P�;�g[>�}�˸b�q}����%m6c���|O�H�J%)��kk׮���W�%9+�l�3�-�Lv��3M6c�\,Z�`p,�^�i� ?���t�v�H{�;���hx)\���h��s�])�':�wB<d��q��gv��n��ͪEK7d�!��\>����	S�׮x�M�1�E���Wo��:;)�w*˿Z�>u���e���-�����s�H�IC��7�卶t�|ˤ��Ҽ�J圵j���nO��S"��.Y��{,W0L�;���>�$�Pޕ�����?��ݪbB�!�]�U|��x�r&&ނ,�z����h\�l"c�Z�b�۳o�:�-I]F�������m0t�( �9�C��e���^|-
�LLx\]^
�62��    IDAT)�~>��[^��ƌ�� 2H=�(� {���3^X��,7�|�?T,�_� cE�)�鱦q���0��Sr�cqn�	 �o.�.�?��<lG2�T;�6~�lG�K�$rn	*�RK��@�cɰ��Nr��^�YI^!˶��$��D���3g�V-�������Oٔ)Sfۜ�l��Y�;��К��\�`�����B���s}��G}�p�Ϛ��$Ç8���L(�{���X�R��Zﳖ�v����k�X�\�*�:��*��3`�J�~�^ms��̦bw|�{���ĩ��-�jq��iם�U=7o�bOo����}�M�b���7ؔIM�L���߿��\��K&:�<�-&D���6�׬�Xɮ���p�&����ʇ����qH�-��ʾ��/����E�B&�it�gܬ�kZ��l�� ]@��a���Y�<��Fk����1���@��X"fK�-�ӧX�B�PO|4�_*�MLZx]�E�� �	��k��?@C*�1�O �!���W�@�<C!z������\<���, �&���/�=���|q(��3��L�c����;��qh
�V�����".�^J5z�b���s}�A�ߡ��XCn�)����e��"2v$�4�<�-�)���騼�WC�
���r�f�2���s�F"d<��Y��L���<��-_��E�]���"�z�s�>������&���?q�,��' ��w�.��?�q��p�)X���m{�^K���>|�r�3 ���í�֟+��`ͮ��7m�y-��؃?}�n���!I�H#,j�~����+����{ð�O8�lz�2{���n�b�Y�h�����K.���B�k��:�&����m�uX�����}�h�
w�x�j��B3��Q3������2���Y|�!��1X̸��h� ���Qy�ᥞqK[��ʃ�M��%����`��R�X��w�p-��%K��i��Z�I$#�?��kf�cyj1�u� �[Dfn��H��ol��'��d|1f	��H.[� ��6xdu��c�d�m��$��.ՖȌe���� �l��N W	d=�U`��9����A�qY8(E���������op�d�K3Ͻ{eT�_����F��T�_�تs�؅���E�Vڂ%묯��|��QD�0�jV3J��	ć�|������
���44��ʜ��	p�k,d�Y ����v���k������w�[�l���h�-���<{��W�kw���nhN�6׮�������<������7�w�g%*p�G�X-��,^do���J9gG:�O���]t�:ˤc�ܼϺ����N5Z{{��,�h{���k/p���!���Sn!/��c1`v����,g^��s	(U��p�O%_��q)�{l_�6;ұכ��h41n���y���	�Ƭ\�[�Ry��5�KU�$����j-�&$�- �1��/n�I���ǳTޅ��#�@��ի�k �xW�?���G��]%�i!����'�!�?5�1t�E�w�=�`_��j��,V|ǘ��e�3 #���^ƍ(%�˼`�S������v;��ɤV)����K��ɂ�x3h�E��;�S*�J�l�������
R�[�\�_�xc �Z������#�g��'/�6�������@E<)��]��kw���v��sl�����������;h;w�l�dk=|�*��}�C��K|�o>c{�����ؕ�Y��)U.����J�~;��a��/�`/\g�B�;��	L��%����n���m��|�*��UW�}�{ߐBCV>3�f�r�X8X>߾�;���HT�� ���p2��|�FI�����юfk��g��#8U.��4Xs�ѡ�/��ր�,/ i�W��(	�[t~BC�09�������H#�?������L� `�2� fx}������E���w˾�U�vޥ�����{}�R�����'s��{?��@/�P �ԩ��`,b�
�]�{M!�
Y4���!�,����ˁNT�<��Py�(���o"^�b��֭;�6]��9�|+����ON�e�W�5�ĳKZ*�`�\�
v�P���'>����V�<ө7����@"��C���K�Ƶ1���b�o�������s�^lS�N����T��d!_��{Z�\IX�^�TR�я��������ܼ�KL(��>��l�o'��e�L�2�>��?�Rq�R���v�7l��U�y��փ^���?�tο����Ÿ�i9f�6]����kM@V�5�U7���7�n��@D�`yPPj��[Ա�57?cm���ԓ�.�(Y�"�Z$i;p��ԓ ����A�|*�'�%Ǌ��U@˟=E#���(����� �����qw>���ƫ�3�/e��r�ԱFh@���>���fl�p�, +`��z����?� �j�����[�@
G��)����˳y��}�f�6@kB�
�#��sqN5p�����4~J�gSc�����V�E�y�ԓ��J-m�M��i�d;���V(�,fiK$�<���ϸR�8������7W������%�Ur��ϝE<�tv���?�|�\k�fl���n8�����\�v��o�x֎w،Y���kǛ���:p��-��8O�����n��m�}���߾�ە�7���皑�>h�����h�_�-�?�j��=��}6�����`_xў�D���l9h�����]w]�����C�#���G��d��gR�s&�{��׹��-�?,(	8�H%���쩧���foW�M'���Ja��	z�v���<hǻ����=���z��8��8QG��:	�"Їw*�s#�`� :�Dy��~���=	EX�H/���*�ޱ�6�S d��R��&���]���O�'�:��O7.���E��wj5�1X$X��s P�]��(s���i�GM�J%cV��_{�'yŬ`U�7$wR�N��K_a�Z��unt�X��ڇ�\�Go��3qy.h x��_�5b)�7�����~N��G�w�0�bǺ�Q[T`qj=�i�]��~���k�`�7\�E�ܺ;��o<'�o�A�?}��n���[N?��r������e$��lX���]�Mv�k_k}�]� h�mmV*Z&s�����~/�0q����W�����V(E���o�;n6�~Ǫ�A�U�� �.#:a���z���E��re����b��sO!1e����b�<��-*b&̛� ��%�p�r�#���)��U����*E��$Y�����g�i8�
t�/�MI� �(�>@�"�o��+I^�Y$��*����0N����2FQ��v�w��E���)�E����N�`'�㆘eh<�c>@��!p^<%��1^��s�Z�	w,Q���Zb�֞c�t�*ł%��n��9e�6s�W�T+�ư�Qǅ�8���˾���9�so�L�ʰ�s�����S�#۰�bPʥ�#v��>��hsj���R%����H5X�T�;�Y2�`�����S�{ىo~�[�ӟ>4��)�v�������t�y$�@�/�\qk捿�z�3w�M�`--{m�Χ�ۭ��{(U�K�Y�m�s-�j�����N��Kd3 x�b�o�8��������@F�dU+<�QGh�^v�*�56em|R��%"���$���Y�N��Q�ki�|2|�zEQ�ꑤ��3��=�p����τ�?��Á?�*�1h��-����1E���0��'��z�� ٗE�W�I��%����3�n���߹�[N�`�(X,%��������@[��)��?�#��8��L���;�4*�2�K
�z;�9�ς���ȅ�&Mj��&{UO/�Xt*��05����T&�4Y���c�]In0���Ɛ����3���:���-���	�f���Rgh\6iG:Z�8���;�����^8C=�����%�^fM�B������/���	���- ���mw�z�WO?���>^ځ�?��^�y筱�_�?��?���zmǎ�]�s��O��d�̚� �R̃��H��%��ÝE����o}k��?�4z����?��?��L&ܠ�����?\�77�k��X�T�$��(Z��)�ʖ�d�>�%�F�^������j�Q����_��M�ZU%�>
62�Ƥ�?������v�n�±������^x?P����{
��E� +@�g�ƍC�d��J`c1�P�*���n���;h#�9 �𦼁<Z����������Ϙq��ba9C�2W 9�sB�: |����I%�CU�t*���>������:}W�%~=.�%K�yrd� �<�RԎ�gt��a��_�eμپ�>��%ܻ!��c�!ཽ���y�HZD=zĽ�'�|��Cpl�˯Y���=w�M�8œL)�����ǝ���t=aQ�$�1�$M
�8���T�/�d��f�&M�	��Z|����n��
�H�����>ॺ8r��ċb03�xXE�_�YX�d��
ϯ���`��m�3��b��~�R����
�Wl�S;�)�b��*D�����$��(�� I�	񏴃�B��`5�� {��6��O@�Z@Ř�l����h�js9o�5�v�\�9- �D�
�R��*�'ޞ�]��Ї>�/Zs>��Cm�c<��p�,
@ �x��P�?�$I�i�H�/c
��j$�
�k�܇J���Ϟ17�}�'qkkk?��1i��?g�$[�p�UJ�fR�P�͛�{����W���L�T�L���.X�Qt-�W�5&Bc�8��x2�B���/�`	�=�1O$��MQ���\�%j<�����$�
100�`WO�3�|X�K���7�s������-�e3Pqu	� {�ej��w:�,2q,fl+��Fݐ��=�)4�*U���X;z&��%����ޡV�];�c��<�Db
@R�/�g�a{��^���>��͎���9O����
p���ͽ��[�'���;T5��0��?���ͻ'Y D��0�G<3���w��|�� 8�� ˛y�1�'��Up�xrP�Gq<��}�W��@P���W�wE�n��ÜQ�"2��:��Mg@s�>G�mBL�RW�y8��k|�6h�Zf�_mF�R�X"��$ǁ���k�lm�Ԭ��B	�Z��嚢��2��_�����Qo�y}��/�o�>扏0���
/H
 ����3\��c`NJA�*�2Hهg�������JMwZ���-������Ƒ�J<�1Ȕ.���dnP&/������->�^kؓ��2�M�'��ŢW�� �%�TUO��F����3+ێg���P*��Y&��~�P���Q/�Lc5���._�$<Y��OF���k��^|X���\7�/W&E�d���y��7������ċ�nx��HOJ�y���&y%t%�_�+�|��R���U�Y'=� 0���1��X�(�THF��J�
Us�1$�Bu�6� |�L�W*��E�%�W}!�����چ,�����β��g�b>��wN���Ujq7�[{�7�
�@������y<^�Q,:<G����s���<&�8���Y��>�яz��W�A�<+B<8�����3��𼠿XP�����d�c�?
F�
�UISJ)%���jG��s*���ZH���AY�|��h�نA�W@�Z�u�	��*�'��Xaox���4�8ٵ;ةZWW���{z:��U:��������w�O�y��b��-^��fϙZ�UF���LV=i�%'T"�\�z�y��' �V�, ȭϺ�������"eч��pT�$8q (G@� c%�L>�ˈ#0�⃪�0��4�G���ƈ
�i�H&�W�.�"���o|�ϋ�EP`9]ŠU��/�|^�W�7��%�CUφlҊyJ�������Z]�>V1yz�O�4�Θ:�/^:y�)�q��>$-66f=��2����н��w�*j')9��j� �澸O����IU�ERυg� .�=F�:��^��H
���P��JӧN��4�z���K@%i#��˲R�h���|��>�C��,��n��i!�K�Ë��L�b�xSVw4�cB�`�H�y���\*�-V+Z__�<�ú�[-�E�@�Ѥ:�e?��a��H����-�g�fOwz(^K�j�s��X5xUp��&`�*�� դ?�e��A����eA,�n�
���$�D�;�� ���Bg����{�2/�`̊Ҕg��\΍�1������,M
����;D���3��x%|8��Ca�V�N^�U=U�٬X����t�rܪ��%bY�5�L�4y�54��L��
%4��~PBC�[Ro<ݛo�Kf�ӷ��Z�0i�'�a���H���ûG����_�Ǭ���L���^f��,m%~1�����j����������#�<|�i�Ղ ��� �@�`��~y���$��!@�Ń�G�n3����眀?n#�q��[�qo�ސa ����Xs�6��h������;CU�\�b� ��ϵ9s�[ie���*�~Z�4�����;��k��P>����C�/�%�幊g,�D����AF��V�!N����ƽ��Z�%ٔU�1D����ǖ�,�EsPF�"���b�x6m�<T�M�ζ
rj���=Q��,OEU=CI��4%ɻ��ϱ��?Ǫ����9�;g�^`����Tz�W�-�V$^���{�*������O9��
������|�	�X�h�U�n�h;C�.�AϙsS�D���/�N����2�O��W���)e��B�W�/\�.^�"��Lhd�������Y˒���-�4�xMx=h�D��;����IKO�[oO������>�S��w����'��b�x谵t�"�3w�U������g�
xVr�5����+��|�O�J>�
���>��{��� HW?��g��ƶ ���q���b�y����U�K��~
��#/�G�D�Z�W�2�D%�k�˜k����Hj29�P=�J)�}NJ:��a���a�ٖL�Ӄ�l�|�*�:s���d�s����H� ��<����3_[�a���}th�s}����
��QZ�1�Ƚ@�To�K�g�g�©F:||���UKގ�������M�z���?EwM���������{��]������ٚm)�R�Bh�iIDEE@D=��S�v��;˝�������"-	M@J	%=�������g~����g��eg7!	p�/^����Oy��y+
/?��4[nHic�nt]j'��Uf5��aM�N9�\@�� w:@l:!k������+�d ��;�c��L˺\�@��ƣ�-EG�Yˮ���?bd�U��D��W�o_��&��q�1P���������\9�����K��AZ�\RH��z�=�G�,;eq�:��\~<֛�#���La�tMi�^���w5�rƿ�y��|7��9�����!˘�ƌ0m�1���H��4Ǝ��c&��D7�`"���L���η.>�hU��c���+ĭ@�����r�����%4�����+��!���z�o�Ĺ���_�O�s���b��kim�����g��_B����
�� �ߵ�\ʙ�d�b^K�T�F͞��c0}���$0��Lw�:y�N��G � `qa�{'�/�+��ͨ�9�#�X�~��e�ǳV"�g=��7n����n��O�lZ/|~�����C7�+��G?F�<�2�Hu�J�R��7o�|��	�.��8q���-��;����m�ē��r���g2�T�Z:t��7�+�c왑6b7�Dp��(�,����� �����u�x���0�F` ��4-2���T�沎���5��w�)�OO���D���`�UW]�g��>����زy�ݻ�ݽ����Ne՘�葿Z'�@0
zy�Aq�V�Z�Jf,��9��Q8ɿ*��/�3�F�Ў����-��M�g�-r�PUgvЏ�3��S1�e:1c���1�D!��.�E�4"V݈��&6�    IDAT1�(+���l�p<��+s�y��i޹RKU����,k��x����R.������P�/5p|�n�zj����+-_�kZ���埓�HDҚ��f��ڠ�!��Kn�~�ݐÆ���m�J�}�D
ȧ�uTU7`��Mx��g���ΰ-]�ʍ�EC)9����R|>��[�v�]mh^��څ�
_��&Rq�T'`nݺ�������E6݁3'�S���O��"/�;}A�
Q�3E44�⤙���u�+M)�ƸX���mZ&�=͖^�[ɋ  *|����O�'�F�P<D��4�!�/�2�����|�L�S����ez	��wU�������_T�qoLA�C��XA��Cy�K�����|%kS�2	���g�ƭV�L��9�I�X�v�Pd�����ӳ�z����,�s�F�P�@߱#?�k�a��V����g��������i��=���'��O�fl�(0��3��"��aX�p+�"
�(3�`+��n$q1K��\�$�:ȏ�y�6V��4o5�SXB` �oni�~p��/���3jk-2oZ�I�B���r��l�
�޹�<_ח�Gn%	 Å�@/K�)������?�ً�h !���2�Y�C����6nي'�z��$Ba���p���1f�XdҎ(�ii,ء�G�
��:}h��v�Џi15*�����ػ7n�?ӧ��I��ǍǉӧXrD8��c*r��,�ٜz��5��+����c�f(ȇ�A��`v����H�6��x ^/^�{����'YR:KTV�>PПn�A����+e�w�V~6.,C�)3%�W1
�L4��*�#)�;p,3RE;��s"{��2�'p�e�_�p�u1�U��#�w��|���j$��رk7�T�Y�R`�Xv�:
�T�hXiL9��<��޹ۇt]lh�c�W?"!Ge�HvPkl���k�oτ@����$��#hjn@.������ѳ�s驝�Rɜ�|(���'];Ѩ#g����`��b?^��!JQ���tv5D�Λ�"W���4�
#p�e����"/i�^
N��i���J[J`e��xj�fJ��o���6y�
�tM�k�tHiJ�R���S)~��?)����N&��N�F�
WYos[�� �H!V"���#hjj���G�豣1��s0bD�-b�&�@G�������7~S`�����%1O�����r�e�oP>eA^��ٜ�1�Ҏn�����|��cu�ً�Q�8sYa[�q�- ���:
� � >�w�gT����}O�K�\b	�D��*{/�����`���x�����N��[
W&�᭭8��3��:�t��+-�i`X6L��u$n�D�P��ތ!	����{L�����a@�]]��gFO�˸ TU$�t�?\L)�"4o�SE:����k�{fΘn)r
R�`��,Z���v�!��"+��O��%�,K�x�����%ȿX阞�;R;��[�>�j��x�K�;�t�"38x��딿�wޏ�+��5��3��Vz�W_w��������RN��}l��4����Ǿ�ml�Ej�|�|i*Ϣާ�x�/���ۘ��|�����t��c<s{�g]�[��7��,�h�z�����wߋb!`����(��DCat'2�j����t�"�[�]��j�c����k��I�����5�� 8��;X<��q���G	���~N����>��!�����b�ݟE^�-�7J��܋L�t�����(䄾�k0m�q�1P�3��}o�ހM^���b-�T������|ģ��r�x}��e�9���(��ln���<�1�&q%���D����5�*�����{����ꫯ�s�������h-��4���f@2�s�������o,J>�6��������]>�t��b3�ѕ��3N�[=�'uD >��7(��u1h�̸#D�~��]3o~`�!��?l�� P(&m3�Ǎ&R1����#9ʡ�;��H#�A��n���Q�,��:�*<O�ŏb!_ dϗ�q���E����X�
pj����ek��Ϗ"��C�_4�y�	���2W�sW���S���Q��A�g��@��5*�2�.�r��vr�}�qN�
�f��h7?n�
șu����}d��d���B
���(�Jb�I
�5k��?]��_˥oz��t_ݟ�{��ʲeϛO���G��$`�u���<�����������u�7p�N�gL���^ U��woL�g��{Nq���8��_@??c�n��P���TWע;���K�3�i�%@K��>AG���5҃��?��������\����p���"��D0����²�F�le�y���	3����)S1|�([l�,�]�|�M
?�{��Pr����j��U%�O~�S��\ ��4P���'ٙ
*�i[���Ի`D~CUHrQ�r���]XR��~_+�+R+�
sA�cˋ�H&�6�Q�E�y f.8���,V/P0.j�N���Q��[��aaN��l��,'��;>��ʆ7��;>�}j����̆�.Y�
l6��X�h�)�%���6z(2�iS�dQ���&P��p�B��}���s��2�>���RiLl1�$`��������i��tPd!R>ւ�|V��/WcB���B1�N�0���=8ͱ�w���~nŜ�)�.�bP���kɕ�ci�X<���_����w�{�:��c	jn�l�*d�7��dZ5}Y�
���W�p̵_��A�We�]����u�x`*~׻�X���	��.{o(&�z ��^���fR���O௩�K9���w���a��عk��SScƏ���3N�~�������sK���O������:�ނy?��;n���,���8G�>��C���LC۲e�|�Q�;���0�����ο�ǉ3Nø�l�R@��G?*7s (35졇�x��i_�U>w�\9�L�,�O�� %�kA{ϯ�a5�8��6H�Ks����ٳվ��B*܆�a����5��!g-n �Ԇ��#	
�S{$�dm�>ט��:�l|SH r��M;��A;߹-r(�]@�.��.�Ի��&
�a�%����	rL�%�����/?r)���!�r-q|d�p,,�C?p0�xe
E
K�E�\|��ˢ�,�Hԏ|��K�_��~��s`��Y9� >Q�	U~���06W�sI:�Ɓ�E&�:�����
~�r�oB�ד
�s~ow������(���|�w�C�	�r-վ�/A!�GkQ�@�W�C��*��Ԟ�P9u�)Fa�����Q�����2�g�����g���n��I�Mwa붍xq�2�]�Y�c-��s�4kƑG���M�X]$���7��'�3}5��_0�����gZ��ITǪp���ٳ�J'��Վ�;6a�ڕ�XҜ%v����ޑDC����ך�g����g�d�YH3�.!���z �+'����ȇ��\���'��``��kj�Vֿ�x���M��9��,�ȣ������hf&����ȕ���g�,ɥ$�1A��1wF �l΁-�P0Rr�el3�	v��c	�sHf҈	�A��	������cڤ ��|�H0T�hx�Q d�����~ݿ$t|�����YՏ*ӈ�'��I�܉hU�	��6|���m�Fb�:��Y��C�e`�-����y}Z]�R�!��v���>��6�����|_�o�~:>G՜-�.����.}���o�G�����/o~(ʆ�xȚ���ۓ��������X�E�l
��*g�����4˂+Q�H����)�bj-���B��/�Ӂ��ͣ���ǐ�¢���g>��F�F��R5Y)Oz�����>S>?���5e>�B.G���ذn��چ*r�\&�5��b���v�L�s�F�Θ�/�+��)=Ͼ���1�����ߏw�o���S�rݼj����$��a4�U�ww�S��d"���6��&����۶�D2�Î])\r�[q�Ygوs�٨�����G$p���[���Z;"�Y ��w���hCie�@�/ ��UN����t����H�ՍƦZD��X~n�u����[�)u�+~�3��O],�@Е�s��s�s��;���Q����(Z��I'�� �pO�����\�֚�F��Ӊd"��a���]�W@�#Lh�K&��8] 4�0���sYz�z���6�;�C�lٺ�R[Z�͔D?���_&ldb<���	�g*�A$\���v�wU�0������%�3�``n!]
9���v���)�ڣ��khmѰ�P������u���;�mn5���F��b$�j�N���o��xI(Ïp��d�w�Ecc���e�0Ǎ�fKZ?���\�,�0v��_ l���xD�Ae%E)�Rp�n�Z?X�_�Ϸ��(��8��5Z4	>7��I'��/����g?kV�R��\<��<r�n��ғ�2��y�F��1���-�͛v"ѝFWg�]~f�<�((�)��寑+d�)B�m�q�n�_�����U_!h��Q�F�s�������v�0��S���ֶ��7�`��lټ�`5V�ۍ�Ǟ��~��f����]�(���G>�[lq�zR(�˿��� >����~��D*gn\o��P�}�9�����|s�<'�e�П�!�u>��[�@�B۷�㩿����{pͻ�j�'���R�r�_je��H����K�੿>�a��8��3Q[C��TbOp)�-L�n����~[6n�I�gb��1�{b_�B���{�X��R˪�d�YhF��T9�aAD����]���>�V��g�Css#�:�4C�
`�8�A:�3Mه4�LWdp�
�x��'�Pi⤣q���/cq(���A��OR� �q[ :;�x�'�Λ;��KY#ΏO!@߹��KMxؐ���������SO��L���5wV�*��P���}x~�Kv��SN��)cM ��a�@�IQ�_)S.��aǮ��랽����X<����8��	���o���;z?,����5F�C���s}�k_���>����Y�ϦM<�^����FMT��ɿ�c�D;���?b��ᨭ�F�Ƶ���0���JᕗW!k@[�5v>�w��^�;v첖�[�mvsPR�z5��_0�{������E��TL8f<>����V�Z�g��N<a��v�؆T�u��ՙD[�&���qL�|<>������I���B!S&ӹ����'�P0����C�Z���Be���J�/]��WҾ��M�.-���@��-"�9�~��Im�\6��/��IG �ڃb.m�j_>l�`A�b�B�y�`;vv��G�!���/��p��@�im�&�F�`�|h2S���kVo�#�=�au�p�[/E>w�}�8�R>f�d���?��#X���q��:�(�3=�{�=��.��L*��}��q\�΋P]4�`UU�4g��JUz�e_۷����?��#G��K�"_ �e-�)�r�&�g9dr��b@�����59n��v�t$��P`��#닙h08ZL�62�B��r���9gOGsK����Dssn�S*��*I>G�y�V�}ϟp�)'cƌL1��ǥ�z}�.5�M!�!��%�-�O<�3�:S���v H� A?_�b*�|ϴ��c��v,Z�8�	��yfS#�Z\����^% � �� +����-1� �����d	�%��#F��v�l��n^��L����-Ƨ����OE��?kּ�'�N�6MMðr�ˮ��AgWk�lB&�N|�����_Cu���.������+ʬ�ڻ�̟!���>Ǖ}��q���o4M�ޭ��Ow��9�M�ݲ��DW��#�Ύ֭k3�߰1�	��7-^��� ��M�� ����ċ;� � ��A�3!�23�߁}��\���Ո�ʄ���_�/�8��Y�8�� ��c<D���M�C0�3�~[�ua�%Ȥ�����Q��ȹwf:�e��4Sr�(׬m�c�=���:̟w1�$KrJ�����ӓF��j<��X�b5��9�?�l�U{�h�tG������,��YtttᲷ���z�I�O*�	�ְ���lX�>�c��/:��=�D�˅�D2�@$
�$�r�0��V<��X�v=��0	g�5��N��R�9b��~?��\���6�����~�aÚpڜ��:�� �RK��y�Ɲ��_1>�c6mڂ����8�sp��Lw�Ͼ/��K��{'��!�z,_�
�?��<�TL;a<ry���A��qə��4��wo
-z��.k=
��rZA�V��>�����Q�>�W�J%�����X)ۇ��~T�W�5�D��/Z[M�a;����wYV��X/�y�[�����N�3@W��5+���s��!d3�\��l ]�Y��E|埾�`�ʺ����?�굫LY�{�/�������@d���#F��|��e\��n��4�8 ����TPƢ����[�+D�qs��x
n��F����n/�2������6,\��x����9g��{�5��m�L+@���[�l���c�+8?�@)n�]���Z�3�8�=g6��X,�7��#�4ͬ�1�7RÆ�Y�ޓ£���T2��_~b�r�����ϥ�Q2߶T+^Y���|��:\�ˬ�]u. O͛�T
�]J��F��ú�m�5�$?}�{}�s'���'�s�JK>C|o����i\z�h���=�����/C6�|�e�h۰�-�*��r��"�NWe�u�.����g�o7���X��q�_�f.�c��|�k�1�KQ�b1��N��f:+5�?���w���0�1�r�-K�.'
�_v�"	 �>֮Y�|��~�N�Z��;����Rx�o�G�2�=�|�
K��h�������cǘ_��DP�G�>�y�|��?Sx���ٓ��E�ބ�e0��;�̨W����װ�����J�+�{*��
��J�KqM�'�?�f�2w�ҥK�eFk��t٩����i����	ذa�~�^�7�����/ K~.�zC�wc��G�c[5����'>���aX�n#~{�-�M���R��b�����A��e �`J�>������z��]x���8rT���]�{M������љ�捛�i��j/����5r�Pkb^��f�?>^y�#l���W��c�a��ٸ��������M �8L�
�-i�}��p���bx��U��3�.�ɓ�@0�u�UV.����o �?ņ�x�ѥ�z�;.B4l��������X�ڳӹ(~0E�P����.A(\�K.��/�p���L��.64<�ebVK��۫�x�_�~�F��'Ok���"M"/�P[_�\&��D���5�"�L��������s�%� VC-�Yg�nT�� ��a�0RE��*{��X���3;����ٵ˄K0A6�<�����ۑ�&QS]o.��x�<�֬^�Y��a��V���teutbյ��l7������*��;���=6�����OPW?��2�v�4����~��]���?`ƌ�s�$:��]�1���z�5$)+��T�a�O��4������ǌBw��(��6!���+�D��h�hG
�0v�N��+���E.�L(�]q_��G�sޥ��@�k�B��ʖ7[HnQ���������R;ŧ�=̿�׮]kץ��Һ�3�O}]�~�>�.��`ێ-�%M7�ջ�CX��{�ص���}�1���Z�v�e����^�=o��/5J3�|>\r�[p�y� �����e�b������2��>�5u���@ۖ����_�N���~��X掸��կb���fR�8����$��1����shp�H�e��.�/ҫ����`��-XH��gҤ1Ȧ]Jlk��6����G�Y��w�!W̠:V��;�X��Id3�u�y�U�H�hEZ��Z1z�K�?�^�;�	�PUU��k���Ï���W]�6�	�|Y�=b�}�Q�ݳq�F�m���mZT8T���[�5k�aΙ�b��#-x�L ��Mhmn�豣-��qs6nX_���~�b��O��@����CJ8A���    IDAT�������l��=;�m�f�X��b�Mx��'��P�K.���_,�b�w��13z��֯{�V�������I�m؄�'LŌ����k���c�����Ƙb�q����B(�@���������a�Y3��\gV�)�5c��񨮪Ǯ]۱e�Z���.�T�~�I1k��Y�`ֵ�y�9��˦����-��=Q��]V���Ą�c�򣻫Ú��6��@g�[�m�Ν��L'	נ=��,B<�,k�ƛS*D�AyU�W���ڂ��H����}����?|_i��!�s�e���[�j�^V��|��!�
N?�t�T�g:�n�Kصs��@���Hg3�ҫ�fV�K/�6���W����܉��.,\�PO�Y���P�oni��������1�A��uj����x�ϓ���ш�n� ���ȫ=��>�4^X��Ip"���>� N�}:&N>U�l����I+A�L�d03D���>6u��0b�H�[�� h@����ޟ\DFJ��~>ܜX�:m�����X��l���w�-s���I��M��L<u�����8ַ����]����)�w�"��_�֋�P��a��5b�䩨�kp�7�70f�<�ϊWV�i�}�jq��������Ǝ3�j��Tr�Y�ʺ��I�i�},��U�0��,;)[�"�ǔ��[u'��\N�֬Ya��-�:;�x聧lc�����\�8��駝�|�o�[ca�%��3O����m�_�����!�O�=Z�����Fw"oEl�\�����+m�؋a��Eذn=fΚ��'M7৛�����8�����b):�v#��Buu=~��[��쬳g�e�0d30�9u��o��@8��ӆ�<i�Z���W�5n���'L7Z�L>�qG���e�3Q�*ڸa-6o]i� �b/,{�=�8�;�\L�t����Ģ�8y*��u.���GWW�7;:��ol.|�l����c�1ۗ�1�_�ֳ��c�o��,)b^k��\KS�Y����T\��ϸ�<�v*�&����F��شq=�a	6mjC!�A�u�˙�Hkw���8��3�٦r�=��w��]�v�ǧ��?����"���l�5uHuw�8���p�EZ��ݝX��9�̙����S�Zpgډ3�3���n�����ؼys��YY���������"�b�Y��O�w���\D��SS؟�}��I*Me����ތ �s�������QG�1�3���N9���
w�옝ǚ�+L㣏���E�6��[�z	jc�( �#F�ńc�������*dy�]���=F����ex������dc˴A�-��`�6ړD%ScGb/���æI�U7�~���u�}�Id#�5���N2_��9f�6+W���V��Dx���gA̿�\��ģ"N:�TD���,hcЕDy��6�>��ۆ����g�Gĳi��@um���#�M�,_�ľ�Фe�K/c�ɳp�qS-B��ة���[���֬{ъ�BA����n�bU8�hh"wL#F�������+���M'���{v�et�btIΜ9�O8��+hI� qԨ#��A�H8�]�����9 ��^Y�Gys,�j2��4Z��q��i���?B.��/����L(�^��>�{v�j���z�`���_��_���Z�5n��3���֯ ��?�9ۧ�����I�?+������bP����n�E*k֬r�D��{��ZP��9s�c���1�-��H$q��oǣ�>�)�Km��A��@�@>��?v�����;�\ǟR*n!�15 ��ј-�Ԁ;w�4ʆ�^z��wS..��'L�����7e���5�QV
NБ/Q!�����ӹZ��)!3��4o��g��|s瞅Y3N,q��L�oji��ˏ��V%�k�V�?����Y�=�l=�HG��Bc�(TU�ώ���S(����c1m7�{���G�Ōf��u����BC�00W���8R(sh߻�,��K^�Ë�9���̓���n��I4Է���,1��Mw�5�hߍ��^k�I@۾5�+��#��3�c?u���kh1����WU��u[����2�}̽�|�9�]{m\he�@2�t�w�EZ��oCw�?��ο�0a�DTW� ��Y�OK�&�
E�2L�d�;en#V���;�c[.�w	F��6�U8X���ᨎ58�K��H,׍ή=�h��K/��SO=m�o޼y���2¶P���Z˰���u�T�,���N��)�w�h۸��c�%f�dShj�Z�2;���YDcUH&��s��3	�}���a�fd�yK�e�?W����wߌ#������Be�y}��3%RhP�E�u��FL�"�Db��(����V�y睇�有h�4�R�o7� �G���R>I���Ltw㩿>a�E,2WR�׸�J������7���OM"��t�3�	J�?�S�֙��,���0�E��1N	ݨ��}��f�o,�Rր5����rQ0����9MEf�9��/e��g���(��L�C�|&n
ˮ�pՕW����@w�����K>Q�.�?�����"���M��M7b��H���e�����;j�Q�2�̾����sK�����_8��0�����d-��M3E.gi�N�8Ͷ�{���m�މ�-Ɨ��O�h�oFu55_f� ��U�1��&�Gx��'��_�����U��,!�\��L��0��-%0_�r���
��w?��O8��Ӎ��2_��1�ч`�u�rM;�&���g?�)V�Y���w-&M9�h�K�D��'��j*(X��	��꘽c&�ړ#F� �l�s�C,,еBM<C-�� 
�<>���z�U��{fO�n�,��9��S���4r��ձ�(���o`��Mx���c��wOյ5�˰��DB��,��*�4���;��o�4Z#�DM(H�z��yy����ތ�5��M��%���ܫ���-���ζ�<���x.����*c��!Z�sΞ��g�RBp�%����?T���1�F��G{�^hB��6���"��ń[r�z�5���T�~��@.�\�}�J��Hu'��@��#�iy��H�B]��n�fA�%K��ɕo^t�ܨ��\X��9������^z)���
�F�lق���[#��G���V�'`k�_����T�.����@�wް����ry\~����>�qJ��aʣ�8�'�p���6[�KKK�}�{1bdS)>�F����N�s��r���x啗��}����y�7o�c�$�u5+����L�|2���p����w[�ͧ?��3
���8��
8*
Z�Jv�>�X˖?�[n��=i|�_G��<�d(�ppEZ�7[�TM����p�w��{�ԩ���>`<F2jst�T�/�\�b������ ���obÆux���o-6	�|_'����	���eEV�`���}�߬0�C� �Zb�V��#���F,G�P$%C�����L%3֓��ʀ廮yg	 E]"��3��T�Θ�
�mNw�܍y�.��g�m��9����UE1˭�.|�_0��B|?Ο���[kwO/�����@� �G�2)OR����`���c	�7\w=�=�XK���c���5��Y�O���B���U[[o�>y�dL�t&M�d������L�,e���|�)l޲�h������
sO��7���6s鳙��L�&��<S�"�*�U'�{���䗮.�<�6,w��=V���=��w��]��f�� �3������q�@�[�8�>��{�\^��3��mWX���9�b�JI�GkJ��|7f8�}p�u�YIw�l��Vk�n�Oƍ�ϲ����o��/�%��s�W}�@��>��������+�.�m��vwZ��EpV���Kˍ�+�̚�B���j�g̜%��	aG����\�Ɍ�p��Ԟ%�պ��b�����������1���q��e���]�������|�Q�Z]���C�z(�'Y���*3o�k��S�rt����OBC6N��Hi�^0�k�87]ݝ��׿n�T�gS�S��"�ý��<^~ �oޗA]���7�lV(Ӻ�}*��r�������q�l>}.�G����ɬu� ��i.g�K�?:W�cj���|�u�p����-U�
�mQ�g��"���MWcN�?��?`Ŋ��;0q�D|�S��2m�iS�I��r�G=L�mj.Ϋ�~��x���ֳ�y�6І��o|Ê\�r:z���p��ӜB�*�a��͂\��R߄J������c�Y����3�\ݻ�F��X����.!��\Ι�Ȕ�}�=����fw��ח����	Ǣ���^承���5�	��ZR%�/p�W��SL���8{�7���\s>yi��p��'�ۇ
�2U*���;�k��`3�>[~WIx����S���]��z���>��h^��Ũ�A��aP�B���O��O��3œn^
5�mR0+�G�}�kMy�0SkC�$כ�޵��$ �����n�����������p�X������<����޻��x9�,��O�Q:���X��O~?��O��SO�F�R���9ܸ�ٕ������fk���ݍ�����J�����GW"� �]�����C�5�����0p!�s�y��>�7�s��Z��2��k�E���6��s��eQ�gq75�)U��[g��q����,S榛n*[w^��2}J\�|>+7�O�Ss��M�Vp���y���l�|^*�&�k��XI��k��(tLP��Ҝ�7�T|f��_ti��#KV��+i��%�3��?�߁������@��>��WZ��?Z����g̭C�g̎���ts�QY���s��ˊ�Kq�
Y�"y�>�?�'&X��N�﷍�~�Cop�?4��c5��4�}ьg�We�X�/�R�����4N��J��1�!^��z\�W_��JD�'�A�K.
�?�;Ǉ���$p]{��S`���ečB<���E4�p"ë4 �ݧ)N���}�ƍ+��qC����H��y�	��ɭ�}n�� �����bޗ�?��,i���:+Ҳ��$���
��j�^W�B�"AR)�J๪ %�����r���T��S�j���eM�	{^�;��	׃,!��[�x��i��)P�Q��?;����˕ƹR�W
��k����ה�s|��x�	k�Ƚa�%>�]�F���ԓf�U~dux��!���h�aY =-��&m�m����F$['9��`�� B��w�X�e!�}��ɟo��?�ϟ`Lp��T�s��I2���N���DN�����G���l�C!z��� ;P7[������U_U�����X�?�~��_ۦ%��%����njC͟�d�,�� .2�ļ����PY�CAI��c���3��4Tj�^�qf��`�K�}��Oa���,��֟���1.fi=��~��aM�XZ���������{���l�e��ɱ&s's�Y��:��)��b�.!�w~�N�JH��Y��_�u�[��������i��X�g8���?�b�0��H>����%U/�MB��� �<=���^ӫ����ͮ�+�Y�\���,t��(��뀚i���$�q�8�Y%*��1��]�a,���{��/~Ѵ4�T��Wr2�-G��[���	qik�*cD�A�=5�z�i�H
��n.��el��.����O�����e9h2t7�閠��?��Σ�e@� F0�Ї>�Oo�Jc��p'��y�FL%Gn����z!�݀�g�u�i<^�Z=�i�󹔦���5ſq�8�|g�>�@�8	2�Ko7��u貚z ^kDs�U<��z���޷T�{��������������$ؗ�X���:�O_2����4.
Uj�	�<N��?hr�?�k�߻�}B��]���]�8��N	�D�f�]�L��ޚ?��c�l+1��tKP�_J�/95p�ɾ�8���ÏW���ڠ��㩽3�[�L#R����I��k��V��S�3�ր����o��4L��ILŀ<0������7O<����]և��g���g�	c+�w�
����TO�+��FA�Ɨ�Qh0���)Gj�{��eE����_��=��y����j�e���d�p�6�;� �  -J�,еT]O���'MS8#�����/,p-y*���#����;��������.kS��ڽ7��w��˔���X  AN��Û�9�f��	��
�)�h��)��{z�!����� <� ����W�}�9�=�I�A	������[np
 �'��&�O�;��;��\��'�+��c$���}	� ��Z��b�6Xa�M���!��@�^�KS�'S>ǅk�V����/�嫴Β�q �+~�ؐ��v����x+��9�Z���)�%O�'!�w�6�h�Z���s ����pK�'ô!�D���+�Sօ6�ib%��-��e�-�|���8-N<���� @@��`/^ %ׁ�&z�M8������;�_�`����C'�D��Sȹ�G����0G�����	D�M
�@�a�����5���xǍ�4i�;�8N�|x�� �%Ùw����j��O�^vdJ�q������'��&L���H�Ф�4���Y�}h�|@#0�4\�+�b�=M|P:�,EU��v�.���T��J�r���6��L-���W�Cg�qo�NU�e�Τ'P3pK�?�2Y��L��1����5}Q�������a�)x�
�x�J��\�C=4C#``�(�}/�v� ���<NBA^�O��z]���zPk��R:����'Y�7ρ�Ţ8�9V� �	�B�-غu;�[�Ě�����M�''�Z�R�zg�ȊP�N�ƿs�9���|��ch��#P)���׊�oJɕ�/OS��3L`�8@a�:��޲�z\�.�Hx1�����r�m����W�]��C{�O7P'�t��'������3&FNYɛ�((Ĭ���>���◿�\r~Om��}s)E�o� �<�N�1���+��Ga�
C#04o�(LռJ�^��8a�8��!y��*Ͻi���1]�B����Ć�ͨ��`/��^{<��J>�P�eeĢ�_��y��s�8[�������	bfN9���햮&>
o~/'�����=�R\4��L�!�#���=�F�Ў �CY@��`vi0�2�|������V�R^�J�
짟~��՛��lP������nG{�#���2诧����_lz-M��7m�|���Y:#'���	��g�2.wJ_�U2��Yy*�~
^�a<��y�����GB7Ѿz��eedV�e:t��������U+ �Y���8�����U�KE��_��f:,DzH'���Xu-�i�4�J#0o���������3�k��Ϩ>����4�]��h����O?�-�6��C���c��)�����z���D�NV�R2쯺�*+���?h�b� ����}R<f�7o�;5~��Z\�P����8�#0P���7
�*������pԘ��
ho߃��_���/�9�$4�c��4u
N�>�N�2X���F&�c��{v��;��U�b����>_|!�?���GG�.lټ+W,C���+״�]��/��a��=hj��_��r�.��S*��6"�<�<I�JA@:���;����Yu$�>��
)�W��C�d���f�J��ߦ����o����ys�	�T��=���d��*b|�ᇍ+I-���,���=�C�,V���z\'������L��p(�DW�v�1i�4�{�\�&�F���� 	#��b��f'����y�e�+��6K�[�p��cxk3�a/�#G�!ѵ;wnF"�i���c��{W'��rؾ'���0>Jb6V�_�B�yK���ok���3 i�#�7}�C�."c%3�xi�io�3�t:C��#vx�W���2�L��� ���q�����yZ���v�a�
;�>NN+z��n�_���N��X�a!��g�KN6�ö�q$ytv�p���4������� V?��R:iI^�7�������s�W�y    IDATq��{�����
�|�tn���s�I�6)������=�شq;
�0�m�c�)s���Et���R N�.R�ra0����[p�h��j����xQD��t�!���n�7�Շ���5+^��N�\�l\3��#ͺ��ץ�;*rO�Y�7��Q9���?���[:gW�<���3��uQ�X�"
�����](ॗס��	�mÉ�N�o�d�ܼu�%�l۲���{�J.�\sK�����m��o������!��z�أ�~���nj[���g�9�|7�n_�L*iڸ?@n�6�����6�cܸ�֞Q��_���)[L�z�[�b@O���"sz��E�����:(�;yq���(��\��o�i����5��`P6�ܲT����O>e��dOe"��(���iՋ?�$}TIHw�S�ߋ���ں6mZ��nrd�ΐD2��ϯB0P�ݻ��|���~�2|�E?��f�Y���D^E���������f{{���}�l�Q��cƖ��W��p�ٳ�Iw`���Hg%��:;��~�&�|�X�������C�`o�(jt��[]T�Ϲe���i���L���RJ�����������P(�����P=�`��hY�1N\<ܣl���6�ai��ʑ���I��fNl]��Mvu�����˟��܃N����jlܸ�{��J��o+WmD6�Ggg;v����/C�%�o��k�������#�Jc��1����4��R�N�~��p֜���Ѷq5�.͓����q�m؂L&�u�:p�)g�{��y���;��'�D3��6w����L�`�L��9*4Sw�����{���{��4������¡r���_��/��]~�=Nk�,����~���]�� ��><f��x|�]�4i4ZZ�a��W�˧��`c�4��+���Ua���5���n�����;�������imn���n�y����������-�i>��`dK3��<^� F�jB�Ѝ�{�!���y}~?��3ؾmv�N`��$\�vK�$�3��\4�.�"q���ӭC�9�	�����;	�n��~�LM>���c��^�(��}�ڱQ��.��7~�������;�q�W�ޥb���g�q����E�̚�`i�3`���]X��"�TPc�捌��G���;;�ص�\x	�=�D�bx��p�-�X:���+e�Z��/ۇk��<A6
a޼K,�3�Ma�m��ٻ{��B��k��<�gG�6lC8ڈ��q�;'��o�TOQ=|�k_3�gF�z2ݓ�AGaB���~`1 /{���6���A�zd�܇�y�ߐ� ,�_���"�̦3�\bꕀPU.��ty��M7�d�B�5l۲{vmEGG;�9�����l�p��֬݀t*�+���ǌ����nK!��������o�����?P�o��#�3a�x��w!	��&���������Ĉ������Z1�ē���	��g������ގ���:�������N�nQ{V������K�ސU���uoٹ����j@��U�C�痦"�h/Į��^'KJǊ�[)�bB��\����MT0���(�v��y������y}��N[��Z�I[Ԇ��[���?�2AҎ�W�H(��TO+D�5��i�0F���K�E(��3a
O�/�@L����;��{Cc�&6�{;�ʚ�R�����uEE�)�j�#�@֬�-���zy8��_����g�{S{ϻ�1��w�m��T\T��I��S3"V�~���<��/�͛6��/����ծ�u*�A8�$S̘q2�u����mہ��zK3�{�R����y��?���R�7��ۀs���ݍk��N\tх��E0�����F�����{�PX���b�'a��3W����R5YuG��6	]=��ԧ,��_�2��f�i�`ж��|Ŭ��������ڜ��`�^���q1�	U`L�`p�L��t}��4����м.c*e8H#���ܔ]t\3���@J B�,��+}O�ϟJ���Ϟ=��*�CA}�(K���^>�hx{[r��#�c����	�us��GY�p��[Q>��_i���t�h<ԉ�?���ΝkkQ���i}�ƍ��̵*^)i�<O���֐�U�\o-���i��IF6Ї�s�g��SO-�K՜j\U��yb�<��wT��~��`��E�G�/�������'5s�?���bʔ)`;L�'A�}�9�=ʣ�c�����D�f�j���{�j�
[�&p�>���KQ_7d#(|����Z��b��c�����h�hR6g)V�lʢ�'N�n�܈�H��,��0�� ��"",��Հs۶mX�x�i��(h+ �����җ�d������Y���H���j=��{��*Ս ��w�۞�@��'P��gg��-p<�
��g�8Â�
��$�%W��o��o6�2��o�G$�]w�mD�e��w�	�����a��s$�x�)���i�eG3��T�Y)ܴ|Ư��e롯���~̸��n�^��nu�i~>�����M���c�# w�R$�2��*�'����-�%�sK�X�I�����2��J�*�4Shm{�y9�V����&��@��~�T 4�R~x-u�b^�O<a>u�[i��`�`�x��kM��t�R�df�=�̳x��l���
�����[��_��_mdAr<�'��'L��"�t⬝R��'.f���/��K+�;�S(�����/�ws<�q}%�_Ҝ�C!ׄ��/���/�	<j�X+��ĤS�=��ng�Z�Ҹz�z�ro�>���M���}C��Y=�<�pT��i��]o��4�ú���4<��;��P�������*�Z
L��XȦM���8�K����c��/8.�P�|�[߲":�6��κ�����y��n���sx��|�,
�����YL,ܡ�ƹ�Vʟ�'���P�'����:Ӧ5!W�c�����'>�ѣ� ݝt�鴍g>Wj���~�,zx12� ��"��&���4�\c}��$׮_��~�����3�
	�a�?�S����Ϳ��q�1��nPo�y_뀱�5ZT�����߼�M�b�}T����*;�DkF��K�Fp_�z��w�'�t*z,� `��:�ݏϨ����;�-�<y2����@��2�@��d&��h���x�������y���*��d�m�w���?�wį���<�M��/���b	���aĈQ&�#W��c�m�b�H\\�r���2k�,�`����	&4��{���{����a ���X��k��|j!��%���9K}-��	[�)]e%u��i����oV��y�j�/^���{���J_ڧ�Ҕ)|9����%
�4�e�!����q�Hx	�5��X 3�.����b4�K^��||^��8j��}w/��9�т��z;Ə��ꪘi�Ŝ�1A�߬�l��N��~�%K���b96����80퐂����y]�?߉���_X�̲�<<_��֯\�\���ϟ���>�ƕ��j>��y���J»�:��B�2d8��I(��k�YY@�5 k�d�RYܡ��^UV�u׾����rl���%v����*� ���SӦ��jL�:3N�i����Z�\�(�
ؽ{�Y�_|˖/�`�Yxp��IH�ߧX,f�[Zo���^6�����W�` l����h;%-?2���}���b�č� 087�|y\�
Ԋ�� C�+]�r��Փ��:s�L+�b�@n-�}�C=4K���"?�Lpj`|~� ��ǟ\���h�`z%�g������ K��UV�5k
��AG�$�;��I��97��xg�mJ����^ם�W�����1�t������T\O�J��}!�PЇ�G�D,Ze׬��3��s���Z�w2�l=���� 	���"1#���lr����u(5>r7�
'6$Rq��Fg/�*�D����1�y�ǖ ���WZyA��N��8����\^|^^��*/[��x���Z��ť�����.Ɯ9s��X������~r�0�DE���U# ˓���pMM-fgry
��)���q�;�]��/ 
�?�p�T_�Kk�����{��_d�h���v6n�w��:l��6`�~̂�a�	|4u��5�F޹���h\,��c0�~UnP��e��dpL����IVgi[�78d�3���M��Lݔ����H3���+�?e-�R��@����~�^KMA`>���	�y�,+l���u��y׊e����r!�{�����5�.���u�}|��<�"Zʱs�Nz|���[��Cw:�T&mY�W�;m��#����!!dq-�)�l�("UQ*~'A�FD;�#���Z�^7��-ŀ�:Ї�?݈��y��'��\^��)6����-�,^�1�Ә�8a�Cʅ�C9�P�"�����82�ɖ�,�8]|ʝ����&L�0wkIY�4�C�_I�/2G��l	���}6�����28_A �w� ~�}9�o�<��XNjE�C�'5f|����P������O��@��p}/_����ƔF#w��@��m�k�C��8�jb�ո�	�x/�W���'���=�Q�,�L��|yms[T����+뽏6�4P��xm���_
Z(���x�Q�o?y}9㓊R������w3Ѐ�(|�XЕL"�ݍ��%BB>�57|F>��G�{��=��Wf�U��?�nP�}Ya��������;�0J���T�Lk��O�TP_{�{}	cY\����|?zo)�^+���|q�r��w���|���:�ڰ���,Θ���w�Wpk���ܰ�C�8>-�XUM)�9�B�Y���ks�u����@n��>���Uޏ_q%߾>��O����j>.�o~�.�\^��b�t�wmmm��HM�	�|z�q�ۥ�b����w>������c�F���8&qӊ�n|����&PB�2���9����
��	��1�j�����	_�ц�������]6P_�� �E#`?	�;ݎ��,A�� ��է2�}��V�[��|pL-1@<��2�4~���ZEWy�5�׼{�Mq�}
��ރ�Y�W�e-����y���t��Zpoփ�8�R�O��SƞR_��y�A���[0�g�xǵ�|�}�������k�k���11��c��w �G�r��R��w����'�&��f���iԇ�k���m����*ȕ4z�p��#����������Q;��W�ل�G �{�B	�$ zP��i7�_6�����{+��9���WC�����aN��{�B���L!fŰBPy��'�Ng|mK�������b�U��S�0���@�����;�C��k����iT����*��c=އ!Ϳ�ٚ�`�/�����^�/W�4x�b�?X
ZQ�C�!�]�J���K�0y}d�݆����}�f=�s�ұ\��E2�EE��"X6Iݜ���S^�}	�y]� �==ǻ�D>�5��o<�~Me��_�����p�L���h{�Y���8��K�;�w�Cm^��R�@~�ײ��!�?����>N���t���b)�3�C� ���>�`	&�B5����|�S!69���A�?�~_�P�˗�*X�0�$ �R�	�S�2�5��e_4����!�?|��/*��}z�?��l���3�K�O#������p.������e�x����W
��J@����A��3o@Ϳ�p9��.�n�G� C����uL_i}"�� P���ؕ�/����^�UX�C����:ʜ�ޚ����3��f���r�i�o�n9�{[O<z>����{�!�<���_(��1��7����qzh�;I�$	 �M)�._7d.Vs*7��+����a��}\@]�CK����+�?}��Z:�?h�>ݩ��;P�t�!�?p�}�a½�z����U1�� ��-����[���om��`��-X���x��*���A��9_�:���W1o��0&�������h
�L.�M��������G#~�@��+Ư"Q7�U���U,���7j(e�0E���������"P�~��������ZB���R�?��q�|t�Z<��*�Qі\i,2�Y6W��Ze����y.�->�ݔ���1�G�����0�^�z-C�S E�9s�(�O�U9����nx�p�d7�錍m&�~P	QV�����|V�6���J�9Q"��p��*k��s<ʬ��b�bU^
�ǎ���X�� �k<�TZSz{+�5��ޞ���Y�益=�{C�Z�'�jo�^Q���G�\�-aV\>_N�渲��\=~ �h����=v�+N̻b�e˞7�qWp6��?��y�"���������q�?W��E.m?F�����zm���>V�=�B!���&-�j`�&K��k�8��*�i���#��?��% T0t8��\�L	�ci���w������n,��R+T��Whv�L�6���U9����K'皙x+O�!is�oW8�tm`iS(�"/���=^��J�������E�+$^���������r�����@��)巪^�hir�Q�H��.9��8q���lh̩�X�TI��
�%�����sz]���~����|g��8�t�QPp���sq�xoS�I��kk]��������)o�s/�'��Ϥ�=�i�ڐ��U��.\GV�۝Fsc�1�2|ذ$Sd�u䆉�k��V�$�[���9\�\M<�p���/��m,G�Jt9���g�y.�{>��r�O:�4nFiuiv_�۷�4C
m i*� "��F!�	���w/�x�B�`��F"�i�RW�~��/�1I�Tۻ��	��	V��x��}P���N�J�7 ���#F�w��W��ss.�R)mb�8���;����x
x�Yc-�d667�S��ל���_ȣ:Ve�.���pu �Q4��
"�c���Y.���������:3-��E�,&	6�#��(���	N	X�{�ݏs�{h�Er�k�;����Ha�߇�E��,-	j��Ƿ��ގ�=^
/��'��s%���g���0�Z���ӊ>aډ�����W�.�h4�ؾ�:s���T�zV�X���q�Q��-�@�ɞ���/����x��>�>$v�3kcU��e�I3��oKS#2���X��Yk�F�-.��ԩS1i���k���.l�B�a.|.n�#�<�ƍ3ӍVB���M$-�C�?�:��~ ��MWGg���h��_<�V�	ۻ����{r3�1������ �U�oV��m�L1	g��ZB��TE@o�W�KSK�Ϳ�CZ��xe�\�Qy���w|G�]���Z���ޝ�_Ȥ��҄=#���]���=w����!��RG����f-!���Xr\ml
���:+a*ˇ���J�)	yZd^b;���8n|w�I�=	��LyǕ�	]�	bY�K�P�{o�Y�)���:֫��~N�:�����~�s����r��9%(�F���q�U{đ�DB�fRض};�y�i�w��Z�Ţ��;|�H{�h�Ŀ�?��'k�h�i n�A����a<�qc�oմ����q��ދ�G����(���c�`˖Mf��������Gy��v2b���nH�L�~�7qQ���<�_c�@n"i�2����5�v�����˟1o�E��H���|�I<��2[%��ߩu^xᅶ���
8R+	@���&�Q�)���x��)�i���8q�]OZ�W�P�}�=�II���^b.�#�l�C�^j���e��r�xP�����;y�P��B-͍��c�8��+7倾�]1�<y�]w݅�/�����F&H��ƙk��#8_����[��yK_x�>�h��D+�q�e��36GlIK^S�7ޗ�p�w�y�)Di�_��O9���J4^��uE�C6���l�Ə,$�}8FrG��ټEc��,Y�[n��L�,�X<F���1a�8�
i��	,~)^Y���&0�!\g��L���3g[G&<��_����j��F^\�7�s���?h��?�'�S�.����w酸���+f�N%�f��xa��,(GL�O-lW{J��s    IDAT��������r�����F�L'����6�}�Y�[��� �!7�c�=f���J�����;�k{�K�5Ea�9�6��K�$���{���\m�����5�\c��X�x�cC3�{��6m�\�*�F�v+-��8y�d�i�r+�Y�.
�qd�1���K�N�/�7�bw,cW,���s����c�<�쬪��N���IH!	%4�]P��2"��"
D�*���S��\D)6H �t, ��i�L&m2s��~������̙3%���'�̜����~������Q���ި a��}6��{�=���FΪ�j�p�~����4Z>��#�;�����f���Bs�8���2^��/Y�T[.ug��Y�|G�\g�64���˵��|3~uS��ڧ��ֲ�Ro��#���4S�Y����9R��q{)��T�E<�|����i�(Bt�y;J��J>�!y�'���u��qo(�\p��Cy�S��?����V��{
��"�3�.���mr��G��%y��X��t��Z	8���e$��� �l�Pe�w�o&��^q��2k��2]��c�� i@���Δ��6Y�r��tw���<��w&,�ΐ�9�<6��p�X�[@�Əf��~�i�%Lb����!|m�r�є�i�����y�W�blsr���qPbl�{u_ɺ1��5`��f7���D�E	��ۢ+��h�ԼV��i��9�����g��5��� �W~�����C�h۠F{�6|(���i9h� �O`�`lX�?��������t���K/��ӧ�����k�W� *��oֱ�/���	L���s�Ygi�l���1�e�*T��9��́�N�lNۏ�X9�kZ��0��DkHU���|�u�i���|��k�T�� �Fu۫~�k�g�ش{�=���|E׽�]�y��=~?��hw{>�=~�}③ll^,�T�������˜#�X�(/��5M�$���u媫>&3g�.�lA�x�or�=�H,��}n};#]��~[2��J�j�O�� ���ڨ�}�r�����r�rI��f-�M�NGd��9��cK}h�������	�S����Р��CM��S���3��r�����8E��̵r���1c�>����#o�q��hO �i{h~F�������K��u�P7���q�  |��6W�k��J1�b�?�^54f�Q������yJ4E��q��&(��Z�v���_j�E����瞳w�/�P��t����E8��Tł������ G�q^�*��;�MPs ���35�ߴ}s�+�Qp�6��)SJ��	_w�y�j��h��Dw���t6�6׀?=|�^0��7ø�m��+��_���9��W���UysچR���i���ӟ�eie�yN�w��Hn�g�zHƍ�˸	�d����U��tN�-]-�\X:�S�����sϒQc��ˋ^����_��͙;��ɶ�+�?�3,�ٻ�&W_�!���ic�<���r�GK>�%MkWIgW�ĢԨ��斤4�k�l6&���d���Ҳ����җ���'�E�hٴ,$۴��'NP�0-�4EӺ�Kܞ��s����cƨ�vb �wM�t�E��pԨ�ȖIH�ײV���h�f�"�\ )���`416\_Z�?�/�B�'�d=�����E��s~��|l�an�]��/��8-LШjh �1�t���CF��o�k��8�]��q2f�o�ͥY<G��9}���ic�o��8KN�~�X���J�w��-��x�W��u{��W��c���uO�ߡ�� ;��{��gk羦&GU�u��O|B��|�+�'#���3F�,}��ڰ'��c����"�iiMI,Q/����$D�I.�ma0{��l���G��?g��&����G��s���#WX"�����By�O�!��-�XA֬]�m1�
��l��.�6�O�F^^�V=�(�B�(,P8bQ$��pL�����Xx�Y4A5����4__s5A��-n�O7��1�	Rv^�����67	b�e���>��kn}�ôG]��xWz�:��1���� b�c�����>����S>���'��ρ%,q�\�:��U>��/�?��aB����� >���O�z�{3Kz{��Ӭu��>�\N#�h�������{�.8}�~��l}A�]q�J�-_��<��{�G�'Ə����)Ţ�ĥ�+/˗5)�l��)�Z;��o�Pԅ��䎟Ȋe�J}�s[�����j�Oz5u�NS��k>.�b^��.��m��c�L�]6nZ+�=�.����d�4��$�y�ؒ��{�E���*~4>�i4`�J�^8M8P�p���;��1���Ȩ��6y{.�j�f��Z�@�`*�8L�y��}��7�EE��iަ���>3���=�����;����Aɿ�	=�,�����ܒ���(�&����k�v.��]���+ 6���o�3��M �
�	�Jc���߿��*�����s�������2����� ������Ϗh(�2���X�PfX(��׭�'{P޲�,i�8ZV�y]2� ?#��lFd�+�K$Z/�YIeC��]'��Uo��fY�b����R�Ap�������i��}��1r��?*�u52nL�,��Sy�>�J����u���ۥ�G�	i� �[��+#k�&��S標�Åޙ?~ɁH��SN9E��Ǎ�R��[nѰP��\t�F[����j��&f,o4�������L0��i���f��`?_�5'���K�F<�}4��9���h����(�Uic��H����l�|6�v�6�c�='��} �4�V�Uc��߿����)��l��������}'�/��y�fY�M���j�f�� ����9��w,,z_��X|��ΎM��ӏ�N�GI"�ի_�Tڕ�A{OO^^|a�D�d���r�ۏ�y��֤?��w/���������3�gvĂ�i�7~��-yU%ڇ�Y��Qrּyr�[����VI&7�����"�0 �➡~��Y׼Q�6o�T:$W|�*}`<�[o�U����׿��=1�h�\r���%�m���.�C��k	_��,zc�x8�/�\��4/_����/[���[>0�Z5�� ��7 �/��|喏��]������<>�җUe��K8�}k������J��ӷ<�}_Y�����6��/��p�z��Z�׵G~��7_�~"��?�|����͊�Ә��@���j����ѾQ2�N��R��C�����BL򹰼��5iK���^";�<SCA~�a���%��T��w��u�=w�}{����/���xC�=ye%�ϓ��T�n��v�X$������MR�Nm���K!�x�N�;�p�m�=�D7�勉ǂ��K������w����%���A9j��x㍚d�S_���y0���Q9�].��V3�r-��r@,�0 ���%`/&tʩ!Ӽ����W�����������2��}��\�3��e�F9��[ff��c����W����TK4�ݗou���r_�9�4}�����$`����Ja��l��K�'���p?����K.��2I��*���חȚ����t9k�#TN$��ttfd�Y��A���@$:.��^eFՎ���77�a�e��Ͽmā�$/�_#k�9�t֙g�	�'�I��Eem�Jy��G�E�4��E���C<DN8�d�0q���&����s>��'1���Q��	���-Ġ_w�u�v]�j˖-�gc��e��+4��6������26g_Ԑi���� �\s���G����1����s�F]�w}�5|����[�3��)��@����?._A(�r��`�mǚ 1N��90������1�[}��h?b�W ����XC�w�;\ߊ��Ӭs�s���WK�K�dlD�� ��<���}�{�+�|��c��j��_�����4�]��� ��g��M�9��s�}$�/j��G{T��կt�`�/pM����M��p����dā�����f���*���k�/��޲�d�i�0�����.kׯ�H$�^���Q�'���x�F�v{�-�76 ��,��,:�a4��{�q�>,6?m~��w�߷LO�2��6�m�j������V�7ЄmL�¡ڵ�|>�����7�-_p�S��P�Y۹lN�D2~8����1�9-⬿5�h�Z���i���ߟ�r���{���)�}�A���5���kв����w��cʬL���a��E5���:���.3w�x$*�|J�I(]�\-�J��<C����Db���勲x�k��L:���Ek)���;�~������)h	�?$17gyW���c�	z�n3R,��ڶ�X��H\6lؤ�(�`8{��q�<c
�>?1�"�.]*].�Ӿc��@o8����w�\����\��U��>ܱ�����w���	Z��\)�u[i>�\>������KHM8p.~�4q��}�9��{Hm]��pF�Ơ�s���W���ߟ����w�a�}/����
`���T؍	r�TzB�ϸ����d�ӴD ��<$.��W˚5k4-�� �Gc8�st!|�ߔw��r�W��C�_��7!�?����0��l���\~��-^~�9c��(�.�n�3���1��3P�ӱX |ƌ�g�$.�x�����߯`mt��[��:;z�V>��#d֮��J��m<�%�)����/��ؼ~�
����:�{�
��Xο��kRa�]c�b�uM@��3g�t��ٔ
2��E ��n�KI7��'�"c��D�|�T���p��iZ������V��b|4���YMPq�JiB���m5���1�n3`����ӸSj�S����Z�T�%�+�}OUU�^@�6|��h9�F���)Sd�3�&Ӓdv�x}�J� l�����ߜ���\�ol�)ٞ��R��{(��n�� ЇM���+�f�?U+�j�HfK�e�=��h��=���t ,�`���{�Z��~D~��ȢE�Jac`���l�d5�,�6����T���lc�{ ��ߎ�7��~f�PoW"���ֱ�O=�TU��A�ɜ��`��?�h��|�8w-��)���}��8��	ܾS�x9��jUϑ��6sa.�9����s�Ľ{ci�����a��s�2~��7��Q>�yv�Z�.b�����'�"ف<d���z�qu���ʬs��E�7i\���6�q��ގ�w�j��MX0C���Z�r������O�'�?��u3�9W�y�1\3 ^vL$���G��� ���w�+�F��?w���d���4<��SIO�>�$�o�]X[X ��kSP���9UM�дa���Z�2�V��pJ>x�AB"Na�},���!}����i�&��~�-.,�-��������������3��g_X2�%l�!��\����J)=y���{���U�H6�@�I8fmb�*KmM�*\q�Ǚ�^��M;�#B��#����xK�=yI%��|>� O{�z�Eh◭T��{�("�|o-u����� ��_ViM���a�QŐ���'�/�o�m�X��p��%�X}|?���E2X�J���p���;f��},`¢x�ꯖ=nܻM��('����5�q���Vp>�f:�v�D��������Wp/��\��B���,��3�4�������8�*�O�n,��F D� ~H�0���F�
���j�Y�u�c��'�.�����c�@����]�\��Ec��p7����#�4ݓ�s�Q?�EE(p,��M��Ꭳ��{�՜&D���1#��}y�m��a�zO)ʡ �bX����tc�z<7֓����	u��w���T�����g�r%,"N�{�iڼ i��^�Z�
7
��7�Is��G��d�?tE���\�4��
��.�;�R��Pi&�����c
"L�N2 ⺨9M\�GhX�
 ^V����
)dz%�����m�2�/+�ZB�{�k����Z�6���4�+>t����Pi)���L^���9��SUU_4�5Kry�21*E���D����x4��H��Hb���9��3���MH�<�Ũz���ϲ��֞�H��	�hB�Ǣa����ϥ�~�K졭g��o�˜�VEV�� yʀ�֥�_�)��o���xn�G�>2���
Ղ2S�d�}��P>4��!3�%�0.	���}O�\�v��sP�G6�W��#!��b��$1�,�6��� �Y�]X�E��D
���F�����-��s���?f�I'�K�w�y������ӱ�5	m��|J��X �>������n2�`&��8Z2y���$�1	�3�tHM�[:�֋d���HݨIR��%��c"9"������ϰ�Q	SS�%ߛ���l�N
Q�LT�y�Q+�ܲ^6nZ��^5-�C���~��d�`��VdN�.�ϱ+�3�����7!�X,��>��-�ʔ9W&ȸ�j���;����p��l�Y��`���9����0]��J�*�|���?�aҥ#��Ϗڒ��*i�L:@��C����a�e2���������g6�.Y�����r��6�Z�v�g�;K�O+8�
y��@�i��o���f��_��u����/
�c)�$ �m� u6��SN9I�<{���Qb##�IL2�uHw�
y��dݚ5���mǾSƌ�(�bA�E<�0�XC �<�
��Diբt��k$'��8I�k$��H1&ɶ6y�OԒ݉�:�Td���/p��̙��YT�$�Ȣ�,�k����O�����DùJ��	'����{�Z.e�s�b��}�����e>=��h��M(���zA�%��{4H�T+.PB��2A����_-��'~�i���k�FMM�F�(؇c[4Y/E�� �B�F���˼���n���P�M�I�Nш��e`<�̢��;��=)��Iy��h�#l��\;�l��Xb���!���*�l��J�G
R�I$�*��:���Ț�Kd����ݍg�����y���6�m��d�*Z�)���J6:^�?C�z���i�I�������vB��'�r�c�� @ȳ:�3�$	�>t�	&@��}[so���$f�(�ǀ�$
�q��aaS�B��������؀0N^��P= /�5��C�R?fQ���2�SJ�?��[]�o�4��YҹZUOʹ�)�ȡ���ۅ[9n������b��L������+�V�i�,Q*%�˨��F]�Z ��S)�ɤU��L�H���t���-5��&"�#t(
Ю	����{�±Z܊��D� �\���I"�"�^p�lްF� O>�Q����G�F���ry=����c�}$"�P��#�$/����-H}�hy�EjE�ui�x�s��{�� {Y�y��2�47'�>3���g�f ��Y�Ͼ�i�n��O"��XY��7�կ�ϱ��@ྍRV��r�Vp�ņr��ou����J#	8��ܵ���c����;��dۇ*�>,>�4��:�ҮA3�#�6���w�}4������
h"h&hZ<L4��1���M|���|�v��U���%�؈�	G$_�jr�Y/�x��82���wu���qN`C�`��c�f=|�J���*d�.���P��:W�}w�"��keڔ�2g��R;a���Tt�`�/�׹�)�~V�DX#��IE�J66Vr����b�F��H��I:�s�x�|U��P�7��8�h�Dv�\Y�4�ӟ������cL�5���&�:�,�����k������?�W�u8���-�����d���RS�ڻ����h�
���~�D\B&�SkE��׈�j�����N4�|XT�pL::�d��3��w��͘Q���1Rp��ާ�|w�,>�i4�%����Oߏ@���Q*��%w�_�K,'s&eD�D��gs8<��Y%C;@�0�H���p����3��)��&��i�f;%�k�����n���52i�$y׻eB�N��I�)��I<�W�@�O\�֑��|1,�P\ґ1��-    IDAT����Lx�d���
jRc��7|O��Z�B��r,�2��G{Qd2
 &<�֦�����G}���e�����G�{${�,n��u�ܹ��'��)K�B�ׯ�iJ�P�����Q=%� ��!��|��r�1����SU1����ē�* ��]J��T{�#��5p'�V�,׏�M���#o{�12��4M��f{4�C��_A('��P(��1��'�����vg��o�|���a����z��|Njh�I�i��pF�|�'`�!�i$'E�hS�lЧ ��n����@ ����,�^�7~�g��F!-�BJŤHO��������2m�t9餹�0e�tt[xja����POH�BB��h�9�	�M�j$����z�>C�߰a��薛�E/�0@�V�۞ c9! �瞫�}ӊx�-&h�ϛ��|� (�ƽX3h
�)��Q�*f{=#��L�(:m��ɹ眧U=�����&�F՗rn ����0�A::����ğ�T����j�/��dD�>��������G+�>x���h������|@b���]'==���+�i�Ji�h�D̳=��Kf�ds$m�f�7�t�.V���o}?���4����[5I�c~=�<��-�J��R���-?Q�?����Ȼ�}ݜ ~�����$���4�����w{�?��X]7��#��vi�u-ᨙ.��%^h�pz�ܿ��Ҳ�I�N�*'�|�����d�]D$L@��7�gP?�����? �/D%��tt�d��[/�P�&|��ٞ��������R�\���@��̔+��s���a�DЖO9�Ufx�[���<s�G��5i�ja�>�VC������k�[	��4t:pN�x��ަ�N3���e���I��J(pN�)@�˚�����YH�ͭ��ZP���=r,����#{��C-r�N�;Zeٲ%���0y��m�=eԘ��Jgg(�L��ؔG�Z.�F4��il�v�=��J����l&/ӧN���u���mw3v��\�T^~�yy�����E�A�%@gƴ�e�}���;Z(���z��'���]�t��g��P<���L^� <m��kl����a��5�7Ż��U	�K����$�RISP�����XM��p��%W�v���I1�)5�#��&��*���Ҳa�����O��:�cͻ0ϡ�4r)� ��>�� Ӝ�I&2�9|#��KǶX,!=]���?��!I�9�a8�>>�E��U�X8"d�J$�O���0��#�=��$�
eb˾cc亥���w;�ʐ�&K�4(,�p�PO4� }�#?��?��pn���_�Ĭ{�@Y�2������n�:�h��y���?��J;�C5�1�M��e��瞑�uM�A��tugd�]f�G-�춇��.��GV�m���9��w�?����B#jf��lZ
��,ym���ҳR(f�.�~�$�HWGJ:;3�����G��
��w��]u�(؄���g��?��j.<0u�i������g�yF��玚��x���P���L$H�l������m������s��(��P�S��Pf���[�e�j����j�)�?�揀��Z�B��֬Dk�P�JN�%������	��p�v�wȝ?��<�ğ�TW����۠% ����I�����wb�)*� D��c�t_����+Y`
ʶ�~�������������}�$Q��c��|���dJA�B�/0�J1�W'k&S����䢋��C�=�~g�)�����ַt�~tc����_�4l�����^��^]$�m%�^'��:I�����#�~�z��݋P��]?W_ k����0i�#2�s��9�J&�?^I�g�y_{����.�fH,"����"�F'��e��l^/==��$��rE�ܒ��%3r��)S�(x[M��i
\�f�Gu�nD��X��K��అl�}�-��K�`J����$�$ �A�
��)���}
P��JZl/��UMG���4v��%����������e'h�������0��|�o!\�"Ų$_�s�ђz�6qٸ~��z�O��?�4�m��e c`n`=����k����g�r�Ъ�<+V�(Պ1+´c�?h�"4��-4gֿi�f���l��QF	��Ϛ5���D׻��V>�����Y�k�>X����(c�D0�P�$��{�{�k_�����8���.�HA���p��4��/�X9�I�tHrs���6˺uM
�(A�C�>���^�^:���K�a�Nz����k�#�}�'ߑ�z���%���l~^�N����5��6�{���v���e��W��#��_$��u�7K�ڍR��,[�^�9��ڸ�M�"�����d�����f8���|�C�/}�K��iM)k�q�8���CY��!��d���z-E��8οv��
��2�k���u�����餝�{�	�L;%Z�,��*���M��NS�?N�'c'L�t7��f���߬\��a�0GaM��b.�%%��d���ʈD��i���G?�%˖J��m�/�P�`�_�������X)�A�Y_����΍ՊF9m�4}ˀj��9�ǚ��?������6 h��Y066�T�S&�	]�N�6V�p^&P̪�s��u�]'+�-�4�cY��%���|�;
�P@|n>����o!-}��2u�x�PN^}�F���¡���s��2v�N�t�j9�'ɻO��x�Ң�jo�,ݻ��_O;���/�s3��,���c"��l��$���r���b�G6�4K{{��c%.�iY�n��sY��]v�uO�n?��M��/|��ݢ�������8�8|>�я
-�xX��o�߰�]�~�W<�ޠ������Z �_5�=�/�w����U6KK���c]���'�3�����e�r�#�|U�'��������t�<3q��)��eu��3;Dy��D]M]��Ʉj�G�K6<J2E���g�f�*��?��Mͮ�S�(7��_�y}[�?y&֏��8��;�	 �~XVn[�&\��� 5����8�aj~��9�� ��bV�YF��=7� �?zf��뚀5*�_��<��g�^��Nj,z�(=�Qj�~�U�Ę�@��n^/O>z���,;�N���AW�?&ٌ��Eˤ�v�4��$u���ǯ�V��FIgw�^kŊ�zn~�����h�l�0�k���CW^!�pQV�\*?�k9��äP��VKWW�s��jd��ViZ�IB�zY�z���!�)g&�5�\SZ�,z{8ַ�
��ޟ$R��8�m�9}�`���s>��� V����5�	p�u���o��匇�EI��֑���
:�!
B-f$�k�Da��3����&�}��ɪ�O�?$!AcZ�?�H�\J���7,�bL���;!���_�1 v��%Z�aS[�UE%t����mƀ&b/Ӝ�Й��|�R�P�7��zt������$8z˜�s����\�	�q� �����H;�()s��}[�:�F�"�L�.9�i�t��gȧ>�)u�ҫ��k�U`��K�B��&�h�x��e��k/���J�<r_i�4V����1���l떥˚%-׷KgwV��m�caٴ�EE�.ݲ_���Vf�h(4�=gϖ�\}�Ĵ�C�����;�y���]�~�jimkQ隈�K��NY�z��r1y}M��e߃T�ǼE�n�Q�>X��ӊS���Ik(���g	/��@7�v�cK�qmAT?����\2W��?�}�� JNi����^�+ڡC�������?�q�u��LN<��D�K������|�.��?~��h4RD"�!j�Nϗ��d%$4 ������}����#	��(1��|G�l��5Do�������M��F� �ti@���}�!��1^>?�uW~,�e�o�I����_�m��˵�"0G��6?�o%�IO��í�i�Ҵ}_0r?8|���<��#�<R-�;�C�.]�S��g�(�����<����̖q�G�kK��K��D��saye�r���ٕ�L6,���:=j�tv���C��0&?:�����n���5�5������~L�j*f����ˡ�'�b��Z�B
���i��M����뫤�#/k��ȱǟ��?���8�j4R1G�q�<,6+&�]w�UJ��}����M��^��m?k:R�R�4.��k`rSBAk�����x�C��崺'��2�
�E��ˠ����Z��K��#WKD���f%�k�p�E��M�o��u�d��i��O��JW� ��GjS�;res���Y<9��\l���%-=��C5�'��W_����/k}�����WU��d���b�ͱ�),�}_\������[Pۦ���%
ڒ�ݞ/�K@���S��,��^������Fa��^��P�,��PV���8� �gs�Z����(k��a��iz]:�h�p8"�]=�|�jIeD6o�:\�8���+�_[.w-�/�5�m6���ܹ��L�]]���]�F�{�{������ukVJwOR�6��\�Gyr�$ź��U�o��Y���רs�ŀ���4v��v�J�{�WZ���A{D`��㎅R��s\s�j�O;.��JN Zd,���u�>���xc�����Ւ��q�:)3D�E���u�jA�l6%�t�$�Ih�g�Hj�<xϝҺa�L�� '��Q�O�.�T�GE����{�i���	z5��aL.2Z
�1Z�!-5"�z�<����_��������C���F�;��sh���r���A�<���a�>5����l�}��6����oK>M��K��l�K֭}U2=mZͶe�&���n�hm]��^�$[���ʵr��W�����p�N~��?�/�KF�%����m��8���m��+���ƙTJ�._���$P��d媥�|��QL*,�t��5������3%��V�1swV$?mq�qN�iF�C��x�%n�E�B�s˜J��ETqkT a�泙��:���db�5;1W�=�5�kj��'%�Z7��U��?�u~��-k��1�[�y��w ���F�eR��vK,��!�l����r��ۥ�y�4L/���4��O��H������<���2�4²q�a)(��B�^r�1*z
1	'F�g�)��w�-���Ev�?�����/�}i��Q@��?��X8u�@���9�9���/��ژ�3�����M��A	%�GK8�q���7ȸ���N)Ƥ�'#>�;��?�s��~��ɫJUϠ�b>���cG�YgΓ�;X�]�m��i���7JG[Ri�P!$�h\�L�*���Qv�6K+C"�)��׿�����x8�}48U� � ���4�����kU��*�O��q����Z0*��%�i�OKWG�߸�E����$	�Õd#;���@�/���S��f.��{�w��х|F����%%�L����_�*�Vj�ƹ�d���E���lZ�ZVZ�IT{���/��/���I12Jr�Z�)F%�-�L^�Q��ǷH"�V�v���b���,D��2F��GI�)�����w�h�믿^�=`N��7�B&5��x,,�L�<��S���OHw��E�g����Ւ��s̱�����3V��^�Q_KJ���������++i�tɱH���0I�s�<y�[���DL��Z6o�H��+V�����HmM��7^r���?�L���ø@�RY$h�˖-�Tp�r%j��vq왃W��ΰ��_� s�r��O>Y#���:"�Y�+�fZ|�UWT�z�5�O�1��<�v8���N�����*g�{��I!��P!-�ѼD�ݒ�l��~�lni��;M���q�$�FK���Dj���ϕF8�5��/Z<>�0��:)D�$NH�>��:���R����)��H��ڧ�2�w��ه~�nԜ�D�QR�`�|nV?�d��Ib�߽�ҋe��	l5��sҶy�,Z���\�R�'64(1z�X]�������=��qB>��_��?w����+*�?tN	�pxf���w�q���{�)��u����%� �ߵ�u��IgSZm�����-�>Rn-��+��� "p�P��/�+�A����í����ꩧ
U�Jt�g�����|�s��д,�?��I�=�y}���~*�%�&M��ft�m⡜�r)I�Ҳ�y�!p���S����K��ه��O5h��<��#T �HB��I���ȑmIm�M�em�j O���Ù�ߡ�7[o{p��c>9����M�+�y����^�����l��o�8�!� ��sl6�ў�T�em�_9.��+��������Sa��1�uw�q����46ޔlO^^	���IM����Ak�\CC�w�}�|��%��C(�鲓��K�_��,~���q�\�߉r �k�]w������H j��3����@�[4�j�A�ᆪq.�K��h��VD�B�}�1b���E�S�`�M�X9�� �j�ѨjN�\A{&S<-��Z^
�n���G�R[C7��� U"q���?Q���$��Ȃ���91�XH�X����G&�W�N)�"�R	�X�n��/�},J�֩	�сo��/L @�@����~s}�].��6N�i�2(��f�TAA�US����fy������N�����r��i���8����HX,��.$+���̓�8q��;Fv�4YƎ'�LQZ[��ҲY6on��x��f|FA�h���O>���illT��駟Bİ
 ( �~�����G/m`n�DS����@�NA��k]i�����s�nL���D#��N1��
��pQ��٣ɴh���ҔF����fc�*�e�xI�Y�G4Ɯ>�Ez�F�bk4^��c��3��(��ZKH��[�C��ܕs{i���\@ohhJ5`�*{��k�.�{([w�y���`_�P�~�����t�"�&V�J�n���"��YY�v��X�\�֮�J���Je8�S.���z'�[�gNc�-���%�4�^�ؚ��"�J@K@� +@`��"���ʩZh��l~��Ԇ�BVl�c�.���`IahF�{ktMY7��(����B���-�6���)�ઍ��E1��r���"EpÚ�[Q���h������x�P�P@e!����I|ύ��U*a�`�--����`q�V��O������'�Y��	|�����Lk-�vMS��������5�<[�4i?1��k�߯Y�ܧi�(Y�� ��Z�~�i����I�$w���to�M��?�>�����̿u]3!���YG+\�a���^T_#�g����Ȏ�N^CE��j�P��ҕ9��<@��tJ�o���n&Ο�Ë��;�s4������Jv��	zr�i�Gi����F� ��Z>����| �WH��m���!� %�+p/}��n��p^.z� 	������%V/ޢN|�|�1XL��s~9 ��FeP�pŅ ���=h$��mnݢ"��Kz,�B.�^B΄{�롅㿢�N�����˪�Z9
n5���z�)���u����_�@m�@f��,q�G�PG�:��h�֢p�X������2��:��]�����ޖ�����ی�i��)�
�1���p1@ӌ� �@���O'Q?<|8?٢p�֤�<�[h^��]��Uz ���瀻W�@_-�-^[&ܠǀ+��ZVV��IT�e-�$z_N������c����7��'�O�:a}�R��i���[-״{��
h�\ֵ�t����,b�Y��+_<�ׅ�|���z_`��û���,�J�P[�(W��qƫ 3kz��a1�~��&J�T�=|���A�?�A9�c��K/U@�o�x8A��"G�h�Czq��r0ƔI���}�`D��@i5�Kt�o�M;���(�JZ�3�\sj��X�l(8@�l67�  O��
�ق��P�[]4�7��0���5|[ݴ�ܒ�\��`ӻ�x	���m�KTSp�����?98�X7Dy����~&����5��E�JQ;[�oL)��>��iHBt�����n��Ÿ�H�p��j���:�4�H    IDAT^6�����2�+�5�K�'9�zDd��b��c�ҺY��j�X�{3��"�'d᳧���Ju�Z}.:���#��t�9x�G��6�6Wt��+; ��`�=[�}|�|;��_�K���7.��V`����n'��3Yՙ��d����fZ�{u�Z��>ڲU[��>�?X�zەuc�����7x'h���m�WI�!ʧwc��p��1�w[��J���T^Vc��%�k��_恵u�ŗh�M>���&	���
�Ma�3a@EJ4U�	pn�QiBd@�Fnf������)��oq/�X�:��t����S���1�����o�� 0��>y��'T`�z��h����"�����E�Q{<C+�`֎�OF��C�I/]��:sQy�·o�c�>[������ι9�l��o��  ���X���p �x����X,�.O?�^~��׭ҡ�c@0��g�}s���������ӁƯ1��a�Q��������"��G���;�('�P��pf������b@�o��
��'��¾l��Y�uiA�Cz����}�l ��?�x	p��d��p֟�S�'%��G������W��͌lo��Qg��4wb�*X 4�D�'���R���_�}�����@@���9��}� v@��G���ZtE��� �~���V� ���<��C=u�IL�s&�h�����O����eԉ/ }��Ea�ꄘ�"8,��L��/��m�;�;�T���
4P�Y̹:,:�D��:�0V;�؂�q�����cJ�O4`ͽ����;�*�"
(� �D����o�� �w`���h����?�.��q5˭��ӈ(p�B5RR���&�O82�o �y-'d8�i`��O�:���&*f��U}���n_����e��$�@���k�6�̀�5��B7�۲�}F@��7��+&<��nA�8G��=VYw�y�Sm���f.�&y��O����������MJ�b�3������a��LR�ke!�>�lQ[g�;�/�7���J����~| >�n�(e�z��Q5��¬%��Q�1��s�å�]t�}�o����}I\  ��唺/�pm���������ș���?�����_3A�s�2<�4�<V5λ�/ � D���0�(+NL: ��z���� ����4\	i���V2
�ǜ�|��?���J�H��!��A�x��O�Sy��ϕ�f����5��R	���uNc�k����RþeW
�E����?т������RN�����Bä�.���-�@i��h�ij7�l�:��6�����@S��z���s�/�dN5{�&�M�0��ie�)�f!kV�m8���n������r�>���pL碆�=���%[�J8A�4����0"�BX
9�/$R��L�Dc	�*/mW��_*'���B?{�y��8.?���8����KNK[8�c��I?���eo6�EI� �|��@ͨ�lxr m�g�]�����a�a�s�lH�9�#HL�<;~�_Z\�{!�s�� �K�,�I��Ϲ�[��3Ӳ`�Ͱ�Z�e���s����d7�d�������{F�1ɦ��Щ5��Q����̿c��y��:Zp�ߪ��¤ɓ.Zpׂ;��q�)Ù��w�6�ؖL~�R�'fN"~])ˠK8 �q��a��ٿ�]�͇fO,���k�+������Y�0�!��6��5Sq[��@c6*��}b�)o}Ѹ�t�d#͔%k6�I(z	S3(KW.%�xL��^��6Q�VsQ4�ׂ89��3ʩ�.kkH�rBݜ{�xUt �͒�*<D���^[� �  �Y�+%Rm|>���-j���c�Um0��/~�EȬ*%�t�Ȕ��B�t��̱���Z'�jWe����Y攥�.��Z�|��֪]�,�r��k?��1A\$�]���ح��+	�\М������`�_�F�;����4�JUOJ�(_t%�'D�g�M�2MC��؝"o�����^�|�K^iO�F��c�Μfl2�M�}5���˂�Xk3K�a��U[�&�q���������E1w��VN<���6�̉d;3RK(�Y��$U�H�X��E�%�l��Tid������u�����й���F�VQ�8�m��Tm�������Ǝ[�!��	�4zh �V�U��������)>����D?B��¬v/}}�=��A�;���>��7�!�W�����#6'��Bm|��9Pko[���y�@��+,�#1a�+f�k�� R��y�{�5#�a� $<��%�Y��VUJ5K8Lq�ٜ�(e�WT.F��?gn?��iܑ+�dS����շ�dRZ���C��8P�O���@��8��^xi�����Z�ro���ݚj��y��dr�jf6��a�Y�C9f8�����gt�J!㣥4!~�	0*�����͇%F�|`!+��uP��Ϡ�@��_*�a����p){[D�k���ԓ�V�֦t\ȅ�moڠ�|0a�٬C^�	E�0%b�V�l��O��F#ڇ2$��n����%�O�ܼ)A?����2����]ˌ�,��?^3�V�����h-۷v/%N?k��9�� ��w�]��{�}���N����K{{��{��e��Œͺ^��TֱA�J��

�]4��;�R�:������ɫH���l*źb�Tr�a�hݝ���S+���,6߲	y�񚄴%;d�UkBR[\��mE��/Eܨ���c�ir�J�/	_ֻ��6����K�υ\�����.W�'�L����3Q*#񀟌�Dr���t�R���|1T��C��Sh�oξ��B=K!���&\��;�Nf��R2�ZD� �q ��0����Yw�%��Y�J��+b/+����/9��O��yC��_�B�q�R\�똓�|ù?C��ZG��w(g���N��\�=�9��bn8�	H�S�_���޴��#��|*<���}�q:��	���K�6.�tZ�@&��g��U~�Qio�T�ɯ5������No�^{[�>9�F�Y,JM<!��V�={7�䒋�e`&�a����SO��5�����{�m#���J6_�g�yFc�-ӏ�/��6������A���~�3uH��+����d��@Y$�Ql�u;�SW�P<�j��#����	Eb��B�I��IM� ��aɤ�$^�L!+�X��c����A��6*�AK���� ��j�J �2g\Oڅ�U�AM�f\Tyd=�X�o%��B��k�s��À������Q�?k���,4r�܉'*��7fv/�`ʧ��	&��#)���.�0�����=k�Z3������_��SOy�~�!:T�m�j��e�/��!3f�R*ߘ*�_������haT�LGt�W5��9�Ǝ-��8]<h_�(U(d���<%�$�6l��-�ƍ3Zv���t�2e�n2f�x}0����I����9I�[����EL5)����~�#��6-�8Zs�j%V9x[V�t���|ø�J#�;^K �0��X��ĊiɈ�:����W��nA*v�[e��骍Ȕ�M���[`�tە�_^x�����'K�~�9Wˆ� �-��X�o�X�<C�A�`=0椯z6}]���A�@�ˢָo�Ws.�{�t���1״y��1׼�s-���<�߫��P�����|ǯ����|��=��x�;$��X,$˖.�GDk9%;�5󺶾Nv�<UN>�4�y�LIC�f���C��o������=�h�3w��$�mWW��!T��#�K.�PR�.)�R�ʫ�ŋ$�s�(�X�����1ǟ$3f�f	���A`a�7Z�O<���{D&P��/��7߬ܧ��i�Cs�����W��j�_߸^&�oP��D���D$+�LR��V��rӍ�	e�x��g�#;7�(�Z�,%����JqMV3�W�O�GKw|�d£�yY�k哟��$�W�����b� �8���"�|筽g4���Eq>�j�6&����9�~���ܿE�Yč�*�;��<{��A�ܱPp�c�0�F��Aik*���D%���+�ʋ/>/�������b�����%��%'�����Y�����mwܮרV�b���<`R��!�/�lJ^[�P�lX�$�74�:^�Ԥ!ʆ��;���TH����j�Z��#�<��$��D�G ` ��Oa��ú�DYT���+,΋���b,Յ�^{P��x^_șF��& #�M�0n�\����œ�	�%&]͵J��"�L�����K.OrRX�4ΓS���h�q��_��Co��~U A��B��;�����l^���~�����߮�0+��
~���`�E�Yh�i�vߦ)݈������ޤ������n�F	0�ǀ�w�o�Է��<��E�*{�֬�t���.��Ȕ����L�SR��e�ڕ�a�:Y�����N('�C[7wʆ��RW;V�zϹ2k������������s���P���&7\<"���̝��d��#�45�����U2��F$��_��^����%��U�WH6�rE�����eg���D��w��o;^{��`q4A� �l(6)�>�Na$:B뀈"��"��h�9�q0��Zp�ݶp9����1OY������Z�F5���)��/I�8zIB����N�����&���ߓ\�[�Ѹ�i<K�M�-�|t�௢�^yu��[��u�����L�Fƕ
�1? ߂{�|p�U-�
��=���QHe����{)�}�yM�X����	���P��Ox��vO&�8�w W��r�a@���57Ա�I��snj#A�|�+_ѐU�a��?�����ʻ�<��?�S���'7���>&���$Y�f���V�p.$�tNV,o�H�N6nL�1ǝ('��?���^��%��O�o���Gn'�*�O�B6'{�>[���5��꒮���}�rһ��b�G�4��Q@���I��KV�l�t."�W�ʁ�5�y��8���Э�;���A3@ۇ�4��6���
Vv�8},�e.���ð�B B���{���-�&�T�B�����w�!����$!�?��$V�h�E��n���}�����eΜy�ӌ�%O��W���ުm~7���.+�ՐK! ��=4C���R�4������]E�WP���]�#6e9	�4���O�X�A�'�0���<M�)ꏡ\[5�2aPm��ތ�7�f�0�i���s�Y��y���/jH)�$���sP�xAa��p�z�ed�����
��M��Ϗ�J��wW�0a�,]�DR=���LQ^Z�D��'JSS�4L�.W_�q�������X����-�����G,��vz�w�ے���+�
��n��U�R��>������C%����HGgR%,}f[6%��i��N��h��<T�z J����}�Ta�nB8By�L`u6��f�F��z�D�+Ui�V�Tw�F�u�Y��EW����� ��8d��xp��J��qh?G����-�~�
�jK�b!,�PN��E� �o�����wϝ'Sg�&Y/%~p���f�'�lU�i����[=k����W�������@ɞ�Qp��E +��h�*�O^�L�[��� ߄C�1V^v�rJ���E�ʩ���R�-�g��k�Q9����?�i�+ <�[Ț����<Z_�җ4ʏ}�g�}�҈�y���SO> ��L�0V�-_,�T���;�e��ՒN�ds[��������F�+������?����YC#��46~;ٞ�XE��Y3f�G���$�QiٸV�ӯ����p8%�ׯ��֍J1Dc5���)�[$����u�2}�n��O~R��L�u�]��ll&�Y͛7O31�������$n�\�b2��-�8�*��9v���{�:�D�X�����X% ���u���)�>+�ʲ(Gq�Z?�A1.���
�;Ϳ��N������Zy��g�ԝgI��;C��5���6�}���F�G��>������9 �hno����`�?XW<����)|+�5j����JM4Z���T�P��}��0�V( v���j�;������w�Y��'��	�TA�Pv��i4�F�S���6�oʔ)�-W�Z"���>��ݥa�hy}�2I�;u.�+J1&���H�^��9�������_�DM��(��?�ח/���✹s��L��/�W���ҢL���|���H<�h8/�T>ho)�es[����ꦉ��=���5�d��Y��SNx�)2w�\��l����'[l$�8�I���eQ���� �-����Dk��PIh$�;��R!�l�тF�M�O}J��7�������DC���v���$�����rىb���-7h=�p�^N��?���:�������k���Y���n!����X5�j�3�ʱh�PD���|�V5�&��	�ٳg��F4~˲-�N�Ž�ڻ��HM�����)(6vߧ�y�{&��V���*�p� >N_,gzPn��n�����3��g?��ww��SO�Fv�e�����U����Q'.AX�.	�H��69���e�Y�HM]��Q�z�J���y2�gräK�ϟ[���__ح����E]S'����-��!5�<���2vLTZ77K&ө��<�I��d�Ƥ�i�,m���+�Y4���n����o����6.)�d�ZV�ղ)����%nX�E�P�j�x��<����(��s^Uƅ	K�x�.��LP��f��a)�sr�)'No���OL�@$=��&�)��o�;o�A����i�g���H�8�Ԟr��^j����4���L��1�޴ȵ�u���/�Ɂ8�yA#P�� �4?+�փ k�5J^
�4� �|fl����~&�����m�������Z�q�o̲���e��ђ�X4��_���g��ǔ��N��%��l�[6�4���O�|(!�6u���kecK����d��p$"x�O�8��t4A�����_����k�q�G�|@ҩN	�Ҳb�bY۴LB����0ц��	��²is�L�eO9������Z�������i�?� ���E��ԤZ6<����M��$y�:O�R_W���7F��DB�r���fiK[�R�Ԍ��lA�����P$�)鍧�K��;S�uǥ�3R���-���;�'�ߩ3f�_2�i��6C�M��<���8uU�7���c�'���"�L���:媫�ڂK�@8�s�_t�E�\�SM3C�T�4p��N@���~�ܔTF�	�ZQ�G��xs����(<p?|�����%|Yة��T�d��l�{����\z?� 7���ɼZ$�|�C���l��j> ��;���
�Y��"�Բ^
���ջ�n�V
��,[�$;M�.�x�I"r�P�k�dR����'Mn�l�]~2�4�j_�,��y���������)�\V�z���<)���	B"�e�<i���]�!���S�5�
����o~�	o���_ %z��g��X���e�Z�5�bc���J��U�I	'�?�X����
�!g*����"!���:[�q%a��J�q�����~����K/���~�kFr����3.��?�W-�j�<��s���*9LK*����os(k�ݾz����o��,[[*��GT��M�lx�>?4dӢx>P`���_�܁�P�cn�u�*`�Z������`%� 0��iԈj>`e̕�c@��8��s�OV =�q^�!�,ɑ��mfB��"֞�� 2V+��t�2hå}l̾���p/���P����?�Q8�n?߳,`��L��1}����Xs+�.�t�GǬ�%^#uu�d�]��#ߪt���O���n��]�j�W���{�����2|��O�E�`�Q�	چ����>��j�(6���n�g8>���+��( �w���i�(����v�M���ok� �C�fX3�j�OooY�h{i��U1/�HDk�G�Š-ڹ�x)��AP����+�B�h��$H�
V��z��,ި�%���K�mG�Ux@��Mڹ�y��k��Dr�r�-�ӌ騂��2}癚<d���9T����0�PL��'>��>	hWW	.��-
�����@��>p�* �mp��    IDATk��&���7��u��h��#���/V��^Z�p����~��G�g����̾"J��s<[ȭ�B�%�k���?�#t�$S.^�Z)+8̧�|�߄)
������gF�|?sl�c|�#�Ep��1��fT	&��a��B�{3G=Y��~�3�j�ܴ����~�z�Eۣ��+��$��3�h����c,^k�d�Z��駟��k��4���� ���4 "X�x��u��jR��BAM�bT˰����G��Z$�m��R@A-�E������\Ahd?�O���_*Gu�V��������z���yN��M��p�$�����&��j/_�g-SX�4,M�"������ |��!��ZrbEdQo��Z�L������7ARm��ל��@?�1��/|A��=L('����� <��K��I�:Q#,��s��!b���D����b>+��wh�}�@����\rnY�����!���uڃD�g�P���<�W���=�����X�p�V���������ϗL^�\��ˊ�tP��zݖk��|Nj�Q-���~�.�K#-�)��`�B8T�����2��U�����S��4���4�7;�w�v��ш�� ��'N{SK�
�lp� �� �X��}H�k�������v��m|f��� �;��wܡֵ�a�<����r�[,,�
͟(����O5�`��Y����f��v��V<�=> � ZWR�Ǭ�� ��������:JKD�]�|�w��P�
�C��a���Ϳ�#���1�����2��Ĳ�X��e�Y�"�3�m��u�^ܯ�c��]q��p���,�j�8�~40�3�@,�El�j������6ܾ�����I����4&?Wt�xE��=�?�գ��}�A���ϣb�?��(�(�or����F�F�� ��@��}~�NZ4UA��������?c6�Ф��*Y�80�o�k�kXn��?B��g�ؗP��?`Z�6��傈�s�'؀�H����&�/��BIq�Z|�%`]�u�����1c�j���B�h>~���a�U:ۻ��������t�Ι;����k'��Y�.6̀��$eaqF�w��O:7���/	���-|�-��P�;X��@�-���>�C�@؄
p�QI�H�����.4w^�܄�����4�j௙����>�8G�>�������i4Ž��{�/�9|����g�h������_\��v��m|�4���t�w*M⃿s�;%��
6͟=�%C�ǣ�C���?�����/ �|&��M���m("�Ц��1v�V� ʤzJIZji�M���ʭ����b)�7�2*��N^#4ο��d{�r���s�ol��i&��AZ9�ɷ0N��i<��o��,�dq�!��ބ["�z���y���8���P�װ[l��4���?�q�h���p�M���������5ZY�h����\+� J�2��?������Qee�.��(h�O�~}Я�����?��1m�/���"�������1`6��2>ބ�Y�������-�������7�Z^6V�5�r�+ױ����ƹ�?jK&/��&�m���<��o��k����w{�v<��Y��%qY�-t~�>�[A��Q��ĩ�B�9�q�.^���M�/Pp_U���}x�,h��q����ڧ+:]��1�o���i�����RS|MD���$�ֈk�u���LR"���3Գ��7�Ǣ}��њɏA��e��r��ڱQ2P��	U���t�6����iS�6�xߺ�Y�$���ri�����m���9�y�ʼ���{�
V�k��_a�̝ss2�~i%�f�BA�0p�T�຦hT���^��_mCb�
̴R]_/y"��!J��x��L��X\2��d�"�0�D�.@�8�[A������ΔS�}���E�@���h��>��{6.n��z��WK(H�y#���'Ml����`��U+��'#�N��f���LHl���3��k��i5�xȤ����󀳼����m�vaw�]��A��A��A4R���&Acbc��I�Q�`��&%	b����ԥ���l�;;����{��s睻s�.;�J��������k�-�9�9Ϳ����!%�kF}�9>�|QHϿj޼�_�I�%����Fm��%�5á�N�ܔ�ɿ}S�?��6fa)Z@בE�@�,I(Q��H��Gs:�cZO�h�,喖���%ʫP*Z�R5�������Th6]��+������V�v�ε���\�/9|�}F@�n���M�(�v��~}Y�M4�a��Z��V��h� �Ƭ�F��|�
���袋<�h;!��C��j+�o&|xV�}h���F�����^� ��x�o4WR:]	{�4ք�s���;�����O@��Xf7��ȹ���6u�5����%�R�m&uX�Z�l.8�� ��p���eZ[lm�z��h�j��?_1�?�2�P�bs:ϱ����8|Pr��ܣ}����O�������<շ��� �������LE7L�?�>ǏF���u���B��{z�����%�ܾLʎ7��	%��Q\X����FC���9��������8�I��;z�	�����J>�s�x��~��i#��8�CŞ���yS�X���T�/4�UOq�\R��l%��$y�����Z�>K�zp	���A��������ߠue|�AAP��R�j�~S'�%��t�3\�
ȎMm�;֚���v `b��5Η�#�#��N4��*�������3.J��b�wliku�u��Ͽ���xĴ�"���hA�s9�3Np���|���M����#m&6�M@<�����,�ac�h�x�����-����I�!L5�#��*��[X5���+Y�J�}�m�����3�i�Bۉ3�8��r�EV��]�_p���C=�?�Xdn���_�MH�(�E��P�f/�'M>�jDT�X׏�n�{������Xo�C����
��cy�0�^�Sۭ�lh���'2��9��4��E���/�����V�o0��t��5{����ҠK�ġV��q���P~G��b�+�k<�(MχD9Gswm-�,^"�Z��ʹ�{6��įJ!�����]��L.���J�5��H�/UҞLv�)'�e�����3�-�"�'����"�������6���o�Ǎ�}���B�KȺ���M]��KqX*����v��I�Xv�B�u�l:���0�XWZ�)�c/�J���8��ⱎq=�SO�	W�Y6h����x���� "���O�6X�B�|5m���D9(�wSP3��뵃^�*;������L	��=ے��׮��]���߽���x�0k�h�T�|�	�ٕW\��>p�.<��q|yv#Գ��R��/�'��M/���2��V|~�p�1�"�?�"cZAʋK�/�����h�$�G�c�����5ݍ�JH`�C2}ϦS��M}�?�y����4��1���=��Ϝ5���o�����O���Ku��\RB�0;@����o�Cʈ���`1�/n4|
�Qȉ�Ʉ�@M@f<�F�?ׄ�)��v��ϲ9�����Vs�fq�fF���Yw�z�����z��{�����Y{�X�O�y��!;��W�UW_bϳِ!\-ZKe����J��s���iU���W�3�c���t.�B�� @A󧄂�q�#s�5������(�&;X��W_I֬(�p�\@�84�,��]2ӳ#l�7�c#�����*����>��@��G-�O�'l�$�������R0�s-�P	<�/`
�#h�0�ͪzVK3g�x���fq��c[[��f"r�
���a�v�y��C\���t�Ig�t3�����͛�l��LUi4 ��>�!|�{��@�j(e]��ߴ������F��JR<�1{�l���7y�>ז���j���3\qՕV*��b�h��p��d�z����r�Q���5=`�r��U�[� �f���v�yo+��V�T����A��0���Wӓm�u��KLOp�ui���5�`�j ��8�\o������̈�\2�4V��I<�l�/�3~��j��b ����<C��#A*��`�
��8��C<�u��h�D�� �)W��#���O<a+W-�r�j-�4�
ax)��G�q�-�jub����}���/*;Sj����zՁ6iR{�$
�ļ�y��/U���@���뮻|�dV�V5o�6<1�h&D� �|��ޡ�?	;���aƳ�Y���Ѵ��n�lB���>��������L��'���כZ ��
Dۭ\��L��J]I3�U�͛>����L�ٝ�ێ����?�a��L���nV�NVP�����~�%�U�g���0vZ߱,v�}�9}6ָ`�r�r���Z����EK�BG&�;{��9^�eŚ��R�8��c^k��q��M�p�Jh���6))8���k�y������B�`��ϴf�ђ,�$`+�'+fvg���=�kE�Դ�JH��q���/����5�b�`}��}r����͜i�����=�2hȿ��/] h�0�u@���c�Q����3�\��뼪'�%,b����Q����k"ph�'�P59�c-��P��Ѿ!�����nSuJ�ͪ�3+�Ղ��^Ye�b�}�Ϲ� M_�ﶓ+#�[�ol	lP�2#�9�����VjٶֿVB�
�$����,�3A."-?��a/J�b��aQd��5>�	篨(�Y�V6�����7	%�1�|	�gǲ+�{Q���9ԭ 1��׼�Zr���������f*c����,C:CK؜�E��O��Z�iߘ����Z�К�9�v~��;}#��}@�6�LV����㏵r�`��m����k��8y�n!���v�񯱝v��
�Р�ʄt��s]��G��u�8���?{�w1��5���as���FĢa'�X8��gu���6�O��]v�e��?Z�g�j�b�r�\��]�Q^e����͟�J���?{ι��n������V��ץIR�: ����.Vi��c.m�1�����V�t!.�\�k]+XB R�&i��˾�}�q(n������jo� ;�}O�q�o\L�Y4�>�o|�y�˦-C~M~�=�Я�_�<�T��ε�Ge��q��N/R���ݾs˷���V�X�q����z��74�R1^��:�����k��bi�2���X��~�z���V����S��p¤�מj��� ������pg0��'�OO,�R�Y 4p�q�<���G�g��g<�����(�+L	�s��$��IH��ў��
GWlֶ�ؿ|���:"O�5W�\����W��o�w�� �v;g��t�s�5���9�T{F�y�����
�l\�5���㙻?�s�*�k��M�Ԍ^ �Ϛ�?���8� @q,���ԱT����:�q��g����}�����}�q�{��l�vKW
�j�2{�
�5����!�r��'Y��SՌ���cg���aͲe��%	���	�1s�w�z�����O>ڧ�����ο��gҡ�+���;���-�.��yOY_��\�Ժ׮��g@�kw�Zg��e,d�]7��;�Y���ַ�A���B�w��S,, �9?��3������cNqS.�)KRB��#�,q�Ҷ8g��CSH�,�m�N����-�	!��R�Z�U�V{-W\g����߸���m�s:q������sd�R2�[Ç�s�HX͍��
�l���_A_������l ���j���O���O�aq7����D8Wt���P����3��~�;q�����?ֱ�p��ҬH��"�d*W���Ъ�O�V�(����~�"5g�;�Ӭ4�o�}kl�����m��.�e�����T���ݽ�v]���~v������6�c�}�;߱_����'�
�fw��9�����!��������v���K=�e*vם��1Gf}�����g\��j�[�.o,���ڲU�v��'�\��ˤ# ���ڦ�zϸ�hw�Ue�}��x�����{*�&֬�����X>��a�Z�)�-�O��uLF[Iy��ʖ�>˖�Y[e�Yq�}���Y���X���l����
�i���Ӹ�뱗�~�ӱ��Ib�{�i~R�:d>�V�}zZ��W>~2>���W��ǳ�F��Haoq��gu���-$���4z
�3�{�����k�j����7�[�����i`�_|ћ��4�a���3�K�=kJ%,xƏ�㾮��2��㿴�P�͜��=;�i[���{�
u��E�ʴ٪�n;�����ϲt��~��Cv�w��@o���hkuBk��tv�SOO�Ɔ�5��*��]��k�=����k��w�f�q���Ru�E�\_\���A[�d��*��pq����������Gc����8X,��;��}�+�WZ8���ŋ�O�bO��9�6u��<E+(tT��4�X+��Q�f �3,��ђ���Gl��휳��JѲ�!K�z����T�Ǿv���S� ��Yi��W�~ɴO<P�ų�ʈiJM������g��d�>���[���O�����'��-�y�3oФ
z�#��z�OIg8t-��3Xԛ#�^�Bk��b��
�_vɥ����}v����4�~��&��k�-�6Qqt\�b�=���۾��bS�L�矟�ډS�ٜ��y�b-ֽv�v�y��򫭭}�[7}�f[�d�V�o�@fϙ���|��������o�\{��Re[�����e��z��}�յ��z{���U����]��?X�EK��+�;������c�|����BF+�ē�'��{�mT6��O⋇��vl4��Q��{���U��P>�=e�4����Wmr[���!K��<�kš>+�)��\K��������v�G$6BbD�n ��,0��|b�Xf�+�v���RSt��h�/��'��3k��o}�7>G�˗��%�?~�����X�ƲҮ��Z;��|�1o����󛥜�����I��}��uk�zT�BTIY�?��}��i�@��g���{�q{��w��G�	��>���Z���Y�X��O����|�������g���]0|��_��_������HMh���9��?��������Nv�uW��t������)'g�L��?����>�����l��%V�v{qI���+݁��ô}���_Kؒ�/���ooG}��s�9�Ezǝ�s�@5��&����n���8&�%�9kC��p�'�(sV��j��բѰڥJx[&kE���]3�y�b��h����I9d#Rd8HkDZ�f7}9O���F&I:��Yk�e�6z4��6�XJ��v�o�.�x�Y�H��͟��3�я~�Aozӛ�W�j�*��>�яz����>����m��=��o큟�eG~�M���-\�B�0��
Q:�b�>���E��)�G>�	�2y�����׾�5���s#譭����sf$����F�O 6k�v����`�-4#)��}ێz��V�5kWY��5.$hX�b�J�^���dE�q䱮ɠ�,\��#~Xtj�ƽ�T� |��g?���{｡v~�����?��c��@�r�nC���%� �8�˰��L��28d9��V��{���� ��A���}�a���w �7��J���d}lrix<�k`ԉ���l#P�(X�P5dU�Ҋ�c�?~z���������� �F�O�s�y��Y�{���_��g��P�(r�]v�;�|?�����O�����U���w��{�lmm-�l����'!�<b�Z���t��s�}�ʫ��z����^�%'�JK��Ϛ1���n��k���'��L�omi���n����暫l�=w7��#�����Qجh]���W�T,�C<��s�z]��YW���~�����;�?��O4��tLS�s��n���������8�R�c�m�m�Qj����Kg���њ��gCW,GR�ӡcX1]���,%�	�䟁2���ޗ0H�x���@'p�c��lL��
(    IDAT�?�K��(IP58}��f���۴i��+�� �i�8^g��e
�D��p�^~�e��>��5�>�����C=�� �����<��`�|������ͯ���cOe=�z��d�
�Z���/��?�Ֆ˶;�t��_�tv��CMY*�<s֌+o����N@����ϤP��M�o��k��%m��?c^��&Y�R�����1�%˺l�=��#�<�@L0Q"�/���F �����O��a2zz�{�v���/Lڗ��I�Q^>!d�V�+��P�V
OQ�7�T&e�T�J��-�.g=s��?)�7raK�'{m�[�v/�:�B]% ������Fxr��(�F��;��ֈ�C�� �G�����-���W�"<�M������W�}~G��-Ͼ�� ����:�i����V�E�����˭l%k�d������)7c��csm�=��O>Ͳ�V��l��η=wH�ӈ�JJ:_uǭ�~e��ء�$y)
I~������ra�Vu-��}�y���?�×�a3��̘1�Nx͉����y�;��mh�Lc���=���k5u�5�M����s��Ga�,.%em�8�-��]8UCMO���:�4 w�d���0%����2�!]	UC�-���U��� Ц`3�x%��Y�>�^����7�w���h�?�n�Z9
�e������{�5׸U���8�������> w�ֶӦ{�t
5����ş�/��gS�~A��;ﴃeR%[��E����l� �@w���[�~�Pr%e���n��ez�m��Lo+:w�\��׿�B�YT�����O�{��n��KG��BU�C>8Ak�Y{G�
�6�3������h��Z<�v�a'g�;&Mqg��������}4�~����JO� m�����;(����3�BMSZ�c�+N�x�>���f�j�rմe�L�R�lE��+�%}z��L�J�@-\tʇۖ�!Z��X����q|�?�S��ڐ��8|�͛WK��8�4���]w��0_(\�3ڇ{�\[;����+.�k�X���G�M��߃F����[
����>$�N�h�\.c˖,�����}�����w�o�Wڱ�g��S���6~�B͠�R3Z�B�����n��扨�&��~g#�'��5�J��\��:�.��"kk%��6���`)0�CC�E��~�Y������MQ�C3!i���������'�͉G�$i�\��@ �s����e�� ;��sN��g��-!]8`d��cx<�f�kc��|��˄0OYX�ކ-��Sx<�����7Y+q�'mN�$И�Q��Q��X��v��w�Ã)ثh�(a8|k�S�u�a�0c�������l�#��Ѓ���q��5�чɞ'a��5�F��cO>�d;�3\9t�X.c==y���m7é�.ϱ��ߙ|#��p�w�(����5���sN����w4mve��7���W��N?�4�o�}|�x�\��0���g?�(����9*�8d�}�;���w�B�D� B��n�{đ�+��	5�N��6!B"u���8�{�>��zp��h�bn��]�A�(�{0�C�q�x���E��C5��y��������|�=
�9߬m�c�B4U(�~��b�ࠏ?�S�[�M���:1YS�t�]p��3N����˗���w�=����/ae��^�����l~�����ӿ̐�s@d@�f�{5ΤP$Q=$xQ�
�5a�� PQ�
�i���%��jqL��S�AN�Ϣ��f���f%��d&�Ae��H	#������R3��I�fB��_��q���7�x�GQ'\?���ˎ;�8��ǧ>�)�&eQ(���I���j�����{͝�WX7�^������K��i��B6��c�?�9��W�P"XZ&?E�H�H�h�7��?�X|�T��k�w�fD��b%�ȐEA��T%�ap���KfS'O���V(B���ڵ���z8w|�����w�?�������0gP:�~�pSwE��3X��@�?ɠ;�s�?ȸ`Q<�����\����, dBs��s:�Н�_Ӑ�I��2�Z�L�6�IP�1���D�9L��E��R������{,�!�����D;xꩧ�+$���U�g3��lsn�|ˎ�4j6�ֈX'�
bwGwRwF�z�IO-�=��r��H�DY:^חe����P�?�u��x�Մ/��!*����N���1|�����M|(� �Bӥ\k�gl�L/��a��R���P��U6�����w� ���W���܅	<K=hk�@�ȳ�?��FB: c�τ��sf���K�O����1���dVk3q\\S�8h8C�I��\ t&�s9����`
@����4:i�ٜ[�ݲ#�<K��Se�e����ޱ&)������� i��ט=�u�{�4O�?���xF���El��'�7 �Eϥ����R);�f�I
�Rb�^�ʞ� 䂕��A\K�B��<#�f��c��N^P?�>��k�P8��b:NV"��t����*�^o�qo	�۪���zgwv�G�'U#�_�Y�˱V���:���L���f�5_���ٛ��f�����X0�zg�y�Kw"pTq�"�bw<�s�[vb͌y��-��ZІw帎��i�zz��@����k��aL�H`p=S���@?J�ñ��艐 H<�8�`�q�(:=��%z�����e�och���I��TEb�h���/A���~'YiB̕�Z��,v�B�� ᭆJ� ����@�q�-��c�T����9�������|��F��+��A����8�J����-���\p����U��9oٲeN� �!�.Ƶ)���q�18�ڪ��,�X��Ġ\oQp��W�Xv-7)A�/kU��h��2؎k����^8S�����?9��e�d, ���N2Syf(�M3�SVl���%tmů����E#�ߟY���3�z�į"!.a,� ?��\����%@�@�1�<�����K44�+bc��j�R�5c�U4�s�����+�����$ˤ�yZ��Fc��i9G|?�7�o 2��<��^d�����Ƶ����t�s���L��?~js�4O=
�+������
����c7��c�����$\{C͸�Wq@��_�[5�O@[��="K�-�t.�P
NU*߃�	n���H�}�e�fp'�[a(���A�j�["��'��MLw���O�_�g�/xA��V�ϱ~�Jh�M�=�;��'�{�ܱf�9k�շ�r�M������9��Λ{��7�Xï�~bs-6W� P���4����z�������2�!��Ŝ�Kۖ[��C��@JA#��M�	L�f���a�|�$J� 䑲�7�.��2�Kg(^�=���@��R&��c�C��P*�|3k�3�y."Ɉ�"�&�l�X)�G�Z����˂�r�eE�;�b���.1:�g2D�T��	�-������U�����������a�$�Q&�%uJ��p�4w)�RP
�R*bZQX bc�Z�VgΚqՄ��sf%�﹬����I�b�I+��%�%�X�/�q}���LҖ:FZ�6�ứ��� ��5�`��e�b�S$[j�{]�Q��1H�;�����k�}��k�����o�|�����p�KQ2^ԣ�40׺�K줓Nr ���?�$3�9AԒ�o��,$� ��K/�ԭ	���.S$���p}�x�l��WG_�E��T YB�d.��2XE��Z=z�(DT�0#�.Z����fB^����ɐ�V�G�Y��=�St�ش�x׎Ώ�0�;j%D86���SF7	�f�w+������6��ɒi%@�F�F҄���8@ I��uo��ב	-gd�o��&�Hi2����^��I0ΓbPԥb�/��͌��o��o\;�j+N~4�v��������!�4.�2 ���_���[n���Ϗ���	'��?�>��>H� u���E� ���p�O�k�B%YƙZ7�?k�+�&�LLKĜ����α�pl�O{q?��P�)����$�>]�L���P��l]W�RI�j���V"O �V[���L����������>�q.�D�
ԳC� ��19��=�QH���o�1標���My�c�&K��)��n�$��H���Ц_AIk,8q�rR�f)��j�~��Ό�ų�ŕ�"��b�������B���ȣ���[G�Gk�}>'A�"f�iA�@Fc���/�Ў?�x��hŃ@��T傡���}��j�r@�0�\�gĪ �\�k�h掁�@�� �i��Z�B�2�����
1�N}��A��k�b�\R�����O�aKD*�%$ejs9B�O[K��9�J�leچf�ҫ�}(�b8�w��>7e=�t����E!庶�:�M��Jоe�H�7��'��ߌ�g�\�M)�C1�|�{r�2��M6�&De���MY4�����G3�5Y:��M��^Z���2XEn�`���_�4�XS��>����$���_�����������?� ^P6��������~F��: ��H�BB|�_p����x�8�K"!��x!<�}xA3Q�W~$i�γG�/��WrO��O �Bk�H 8��K�-Yh��͍Rj43��y����'0K!n�+�)�y��J�`�,��RVJ����)���Vk�%m���-�
���rnsC�s���hj�Y�(D��f�'�\&`a��Λ�=��7���1��] /
��/N��z �OR\[�!phf�5���~΂���#-8������^,t M\&�g�ӟ�4l����e�������C�w�ԃ�'�ZOh�O>������
��K�U���hd�}������՟�ٟ�` �n?�n�kB��~���=a�5�r��w������G<;U.���K�q�G��1���=��8���m��b���L�c!�fU�y��UI�80���2N	��%�[�q��L%k-�i+W
V�!KUKVv�?g�
I ��M��$�������]{�uȍDM)@@J�h�P�"D
���w�ڷ͒�"���?g�PO9[Ўpx[�qlB"7(� x��is0DV��c#��2ɘ�\�SE��h��=�G�}��~#���黥5YL�hƸP헱!����g,�k�Y���a��)����:��g� ܧ�z��J�_�0������q,V�b_�tVׄʁRB�#נ�V�@2�9�nR�@<� E�i��\-���W���شO=�C�S>p�Y|���U�k�Vm��w�=����V�B�bm�f��Y;%*I�*K�:�g��a�w(/���=g]��XO����2��;d�y�1+.�D  8?q��2va��M�3�q�C���O�	�GYh���~�8�B���0���L��Ϙ9�	�̥Y��(&II4H_6ٹ�ז� Px�����pP��<��.���¡x�E�L#8�-�x˄	�F���_^�/�;�28cΟ���
\��g�6�r�\1��5'�Ua3�����%*ǠBݯT� ��b�E5ȹ����|�r*� �i���7���Z�f�U���Z��O;��8�Dˤ����Ҷ�������3@\�;��mP'h�:q�А�,S����u����ڊ]�կ�j]+��Zmw�'§�D�T�X����Ж����c�r	氖���'�x�+�̹B`����Q؍a(��1}�hMh�oV�G`��
��s�:�N8�P��2���n�ZK���|�,��utLu��{���2��Ln3�̖>���駟��R, w��WOc�_�U�P��Sc/�L �����e,�{�t��
�Sē@_}�.�Q\��=�� 8K��zNC&�8BD��d�i�şK�������_�Z�c[��5�nf2U˦�V.��i'c�{�IV*�[*M�i�Ǟ���@��5�O��Rٜ�R-6T*�50�+�T�h�){��Y��+�h����k��?��m�]��J�^�)�9��4�VHyd�Lr<�p�y	N�W��?����;��k�S�T�U�,m�&4�7��$��*!��s;��o��P�![�b�����قE�\.��D�;��C�SN���lk�v�B��tcΎM$�_�_ٿ΅��A��sbPP�q3���P>g�vz��{�s���|�Z�W��}B��?�K
@����]*�������6�4j�6'?���:�F/͚��lTzAsͺ��(�4u�g���/����@kF��^ti���(�_�g$� A"Kgx�|=#�'h��n �{���٩'m�j?�>���l�v���<CJ�t��Z�m��1�Z�H-�ݷ��Y�n��"�m��Gm�o��RC�*g���h���w,ߛ���Z��=���J���-Mt���[�i�C��d���Bi��j�+�B����ʷ_a���a��y��.��ϡ�at����;V`�����#�w�Cה�P��'4�7��_�(��g߽�?��&Mn��U�����Gg��5�kQ1LJ�[�v��Î��:�'��&�0>%6q<�t��ALv'-��@m&mQ��EM!d����أ'�V:p�4,�x����	��T��c	2�
���" �!�/@�˺�8]WB�ϤM*�?��ba�k5��e��Z��H8�&�6���&`��1#��!�3�ϡ�U���~�s�k�ԓ^m�r�����mmڶ;��`ي��M���e�mV,T����1c�M������P���gh͵Y��gK�κ�.�j��ҩ�u��ؗo����X�rV&��7��g���X�g<'�G�[Y� �A�-`]��>�(��u�㼟5c;kɘ�p|rr�Z���Ckٌm��L{͉����z�C_p��9Y��Yi�����|���F�>���ʦ�6{��v�i����=��k���^m^x�z{{<b�D��F*e�Ww���C6u���_��ӎ	��~DgP���#D���	Ĺ��o~�I8����I�
����ϕ���S+������|ST�P��w�ѵ��w��a`�������@1S8fY��.Y /�'*�*�����
J�=�/��"
(~6	.�d�����xw���NT��e3��}�k����J��*Ռ��v�Y;�DҥlҤ)�΄օ8|{{��\�����v�P �{lh�ZrE�Z1���4�c)k��]f7}�[��b�T�U2P��T! 4t��=6��Y/�5�
�V^���}���3J�J�s�8�^RV���.[��{�鹶�7�t�?T,��@�֮[o�춧�~���ʹm=��[o�x XF�O'y��}b�z6�͔I���iӷ��2���w�=��+v�R��-z��}\S��ށA�Z�e�r�-�׽�ӳ5�8���-��ވ� �����pCy�������/x���!�|,ir,����j�c���Oc.���{hl>i��$��<v�BH���c*�O�P�S�0�"�!v��z�N��K� �yLO�7�*�/��{Z���;#g�$�3���<�4E�o�R�>{����I�=���>�fZ�c�^��nX[K��������R��P���´��&O�/�io)YO�E��/5+�[&�f+��K7�a��a��"�ԁ��y�u�A	c\Q���%������2��>����m�f�>�kKY�e�[�x�w9�500d�m�mɒ����V�Yo�\v�t�V,V����[n���h���&4�7��K�1lםw������X�w3�?�y����c\SX�|�5Pu�?���/\l}�f�W��~�b�z׻  z���Hh�LL6� �٘�9��u�U�\킀�!�nEn����8uƂ���?6�v��f�c�޹��6�w�99J�Ҧ 8�x��f��`9�b�&���u�����t��9c���Ɗ�QB1m#��A4�^]�T+���X�H�q�;�3�v�%{%Zt-����
���N������'a�r�U���.Gٔmw���oZ��B�J���th(OC����X�0��{��Y����׻�o�d+���7�ak֕\�SF�	�    IDAT�����_�>ߓg`�E0�\�`�PY�ˏ�dt3�(x0X�KϷ_?��}�����Y��s�u�;x��l�=�س��vؚ�}�������v�k�+W��<�ŋzm��"�W���s���lOw��F���Z.�>{�e�|�u�Mm�������c�y�ў��l�"����	�d�֓�%K�Y��j������~�����v !�����y����L����H<�y��>��x�v0�C�9��scC��[��r�4"J�F��{��>��̝�hb*@�W�t2_
	i�Ҩ9^��|��/��:�,��U��}E=��~=��Gk��R%(�N��_^1=U�p+%IЮ��Y �h�T�:�9�N<�(�z�Tm�=�:�Z�gY��/:��	`$w��������� ��YOOޓq�����Ֆ�-�j���{�k߸��v��b��MLmE�RԍVI<���d=u�Q��o��6/����C^y�^}�}��f�n%�Ս"8�����_�mGq�M�:ٞa��*EwDS�(��g/.Xj��$[ݵ�֬�O��=J�ZM���{���|<�-�a%`��o������c{���X.]�%K_�_��#;����R�ŋ�@G�˶8߿h���ڳ/���~�Wgd�����?\�h��ꪫ<��+�q~��pΟ"]J�  �(�J�l���q�V��ǠG4�Nr��$��o�� �l$H�o,�w�e����˚a��S�� ]O���|�)��m��@�?q�|VuZ��)�ɲ��� _����	�RB���[b!��#�w���W!�
��5�,U7�v��N�לp��J�VI����l��if���0�=X�sV����RgK�����2x����P/��
C�V�H\%m˖���[�ۖ-ﮁ����o�F�����b���_�c��O~��W�r8�x���|�#���z �������~�=;�l���J�h�\������-���Yת^�d��>�i++V)��ӟ��-\�|�*���X9���\�p�V1C�Y3���|��V)z&�7�q�w����UK�o}o����D^�p��*-�pi�~�1^G�����(�t��l6x`�Wac����Ss�=6��Hӓ8h۪�7����? ��;@2wp�l�_��מm)�Z!���UV��b����/�ιd��X����,rBD������B8��X��Q X[��v�\��ƽ�YOj��#Z��F����G���R��R�;o�T�,�1�Q��]��l������9�
C��ɶ۔�{Y*=9������\�t�ޝ���{�X9+���0���a�������
�P�ǭ��B��5��ׇ�|Ya����{��w�XSO	
������^W��f�c��"�W�Xh���ǎ�Î3l��'j��Ht˶�ܧ�Y�J��m��N�go�¦M�i]]��N^�腭��h
�L�J��I�f�d��Km��w��\������Ͼ{�`��]���4����x�R��Zo��%{Ӆou�`C0�ԭQ�8����cs:/�¹3��h��).��7��V�o��f�% H7��T�C=T�×FkYr�rGE�����
@0 ZD�!���zj�E`��gb>w�K�)�A�?k�{B'��  ��L���r"J@�kp�]w���p-��~yQ/�u�f+�(4{ u�_JX������W*���%����jf��b���#Z����ed)���@��U���r[�R��[*I����c�D�� 0N15w�Eفh�W嵳P ?����R���B́�&��ŖIlĽk�&������18:�l��նx�*��ڜ�7�QGo�t��>���緿S��}��U=u�J�&��3O�׿�4*���}���l�e���L*k�\���Zg+��m���|��j-����"�ŵN9���j��{�q��a�c�N��x��s����#(-Sa�lZJ{ �R!�����<�N�����bߍ��f��W	��:�ی ��Z9�ro9��q��g���# }��|�߬)�G�>פ�3k�sE��i+�D�EMd\�H��C�C�1]�G�����p�|�G+/�<>�R��M����J���H����B�E%�s ��f�3BI��uPM	�I"��$y�9GFio��G�n���<R�A@q����q�E�\��o�r+��.�[e�kW���-זAY�5k�=}�1y���^o]��-��oo~�%�݌�\J��w|�~����5Дc���������[�\�?�r������9�_����6�×����O�`���ˎv��o��ӦX�2d��=��Þ���i���l۩����w��;ʆ
%��@3d�C�F0��DBew٤�+N��墕�!���G����?����3��(hȊ�Q��;�K\U1���#iD1���hq��@������ơ m�K���h��%A=)	`�U�
�qM�����x�y���`�p" ��{�zR���� �zQ#	3W�+������'Y���ݳ5*��y�н�
hᐸ݆'
�L% �?k�U:C�^A�'1ܴ%� �u��ט�g}0�c,E�$OB�����c0�(x�;��x㍶��)�^�d�-x�9[�b���-ז�l*k�C�6y�6��:�;�H���N��jU��t�Ͷj�jǯ���`fwv~3ߓk�hB7����N���>�.��ki�X�z+�����'6�U�8x�A�ٱ��i礡�~;X�s���J�\B����4O{�����'_G�� [���S�WR�X�������U2��#�H��[���}x`�`�5��.?�/-PU,9� �@q,稜8�����Y[�8��(%\+Dk��*��{��f]J J���)��
urj��֨k�������Oi0�.Y�5���(Y����ܡ����h֠Jl]���U16�����7�D��+�(g�X� ���1���1c�Q
����lp`��Lj�+���w�e�}yW��:m��6u�t;���m�]����^f��q������En�F�?g��������S0C%�8��'���:�u6���z{�[kKp�6X6ko�_�Y_���P��~�;U�A�x*��BaC�,��niܿ�6�2/�H�M [��9�3�w�^�:Ná�V*��ŝ˪�󷦕FmE��7���}� �F�����UF'Bց�����u���@����7@3�:rfs�"~���q>���ǰ�P�$X}���.r�A.��i��qkP��AH{�ɰu�ţ����M\���o�;�� �[7RR�sr���Wj�FM�4X&��J�HI���t	�ׇ~�)�%@��B@��(��ߡ�O?�u64H�G�r-T~�vE��E��nc;ﴫ
���p�i�{��ahO�I[�H�k�WR�ab�>�;;���ɿ��.6}�v�h�y�v�i'������!U�g" 6�SO=�� ~O?O��)ڇ��?�����W�£X@d������
4I( 4:O|�V����<q��`ߏ��=+�s3�6���%�� ��ﰒ�S�$��|B �D�p/�s� 7���zA0�9��>` �1ψf	�@ @'r,4��s��\�Ǳ�[օ ]��m�X�xP2�څʀ�E&?	��9�j�2��ƥ��$�zR8w����	�>��B�}���������哀���� M���>hN!!,K�qf?3�8��8�o�� 3?*���>��{��z<(ԛ��z�ɧ���g;�8��|̳��|���}�1i�Sy��|�������Γpk�ʷ�C�'K18�B�謥� Tڴ�^g������Kd{xm�G����9�=�����#:�J�|1� <�lhLB6�/���������9�n��?�(ʹ*�K�s42�wM�R��ߥS��U`���%��a�3�̭Z�1�k����3� ���h�h�QQ�P�3����7�FP��$�?��5���M&J���V3��Ij��+!�)���q\g��c�<)����M��Ki��s�GO�I9�c9��4�kS�f��u��(��o��M4��$%�k��օ�O~��v�]w�~���+Y�{V����gM�A	P>�"�v�q{;��cm���9�-%�2tt��=��S^.~ͺ���*�vL	��dF7��gΚq���~S�q��s�t~�'��htͿ���R��b�r�!�'�=��͂$n�P�+�8������C(�����a���� �Kj7�=4�K.�������%{lb*�[aS�V�{�D�H&|�xw����"`�?��^�Xjr�h���������@փB|�+*��կU{L;q�k���N"����*�W�e���RX$|�'X<	�'�S��寪Y9��y�������0�k�W��^�`��0��2ou|-��F-�3�{l%�<f��|�U"�'^'�k2uk"~�v��; ��׾֕;4*��ЩJjd vS*>�
��P<4���|~�uw��|�$	��o�R[[(3aqo�Q�����C�XXmI|�����n�9fk�xQq��c�ɇ2@�3���dx>��N]s�5�9�}��j��7׊�!XDlLg@��������29�1�[m��ix��f�% d�|�S�rK�Yw�$?%�c��p��E}��qȋ�q�^��ω鎀�8�Ѓ!�������6�~|l
��>r�J��X��1��V��յ�@��f>��H�c�%��أ�:�kn!9�%P`В#�?���<QK�a��k�BeCoK�w�]F]\�}��KC�N���t������S�=����'���E�/�G�F��<jxѲs�׆j��˨�<��4�S �w欙WOH�������{.l���}#0LƆQ	A�	�b�VE|8Y�4�V$��=I��?�s/��v�2��Фah��Ѧ�
8��B;}���~����}�V�lGi����Р�0Nd�G[4��� x6At��8�3��˓���Q��J�s���$F��s��Xq�����߯��$�����f���b�������D��3vs.kF��a�0��^z|N�L�� �5Ф���y,(�^@>^�̔�4p�Ԭ�@Ŗ����)f��P�m���9�=��W���$5�j͉�1V@��/��-��ZK�
�|L��~�(���u�?�/��{Ml���%ߓSc�	>��l��R5�lD�Ol���i�M�?N36p~,���ȩ��� G�L{q����Eb
a���"�t4&(�[��-�������8xd�5Z�5z	E���B>c#�̜�<p�18�2!��)�'�G��<v��3L~��㇫e>��蚪���̋gB� (P�����<�� ��j��<E����B�9�lt*jJI�y��x&	]Yc���"�D=%eFV!�s�@"`�.���l�40��1|ox��Эk<�Ϲr�K�I�3ỏ,(~���o�A c��FBIyc��U�c|f��	���,�$�����w�ynRKsd���]M��9*-K� O�F��C{h�j�)Z��Y����{�:�+j���F}��^2�"P�[���E��O�<�|U"�K��><�B$�k��]V  �s���K��gNI(㧴a���9����"�T:��	8@�8��?I�=q�a"���z�B�)K��~�[���Nn��-�z%×h~P���Pn4�MDՉ�A`IS��r�+p��\�����O���Xh.CUP�:��Q*&�w5=���i7����+ƞ��	sc����x���6���k��fb�'0�"U��T��C�Ģ�糁y����)h]C�����1l�Z�i"h��67��Xm�,
QͿV#q��Y]�.�q/�+ A�:cD������.���g^T�pt�o6�cO/�7O�J�:J�����	o���d����Љ����Wq�����6�����B��f��y.��uyv :�s�.��_~i�Ϻ�'M�x�y��K�9�Mx�����j���P~g��x.��b�C�I�"��zI�F*ž��y����8]��>ße��Ev�-��s��4��p�&���ԯ����#+T4m}C�F����'�7���Fm��i�	���8�e����E68P�����j�-Pa�0@4%�H��8�
w��y�������/oX�Ζ�����$����d��Ҥ���pH����qrj��\[N]�<7��	ϕ0�W�) �f̵ J��$.Yrr��LkO݋��YJ�R�g	<���@�����}xO<;�������d�] �:Áy�A����ȓ�@�B�q.�o�w�8i�|/�Cd2š�Z�::s�G��"p��-�_*�C���}�(����3O�z\���W�%���4N
`.D5SNF 
5�^�~�
�1���wD��(�A����h�A&���K�!h�ld5��si�V��1��,l4=ř�@���V્΢��rP�D�/�7�m��N�F��ܺ�k��ъ����_��X����c��>�y�<�( �U�8D��&����̭曹��&�Gh�P9
��oU�Dx ᙹ'�����e��s:R*��15%+�u���R3���|b��L3�C��,7�A�<����^�7[�zUT	7D�[ �Q#Ifq�ŦM�nm�>��W��/��^*ݩ<��o��/�#���=}&z/����b!!�b�<c,0�	�f�~Bk�c��7�z]C)[� �5��Y��@�4|i��6��r�rY ǰ��81�R{��K� &��.�f�� ���t�fZ�,�!@	s>�	����|��4n�A�.m�EEc^x�>
I߇����?~�[J����o t�K������;2����X����,XB�S�>�g�����EY(�RJ �
�s�hA�N��O����`=���f���F�'` I�c>�`��#T�>=!�*�)8��Җ��l֬�m�?�Ψ����CJ0�D���t�8�'"�_B_�@���W�ޯ��	��[���sD���#��3g͸rb�z6)�6q��e-�ZN�@ҦT����X�\O{�簨��T�M���a6�;��@1�2'��M!}'͟��YX�i���኱�"EkH��Oir���U$��;]W�%�CTB�T�ȱ�N\�8%����Xm"}���T=�EK��E;4N\Ka|�uUs߿��Dhh��H�_Y�������xZ���3�|�s���y�=.��g ;B*	���yF5o��ǪDH�"+ �
���!�<3>�I���M��g��)�Ce�1��\b��GF,%O��޽��U��Ο}Ʋ�S4��a�n�������-_��È��?/�j*��p��֐�{	I	,�X�|m$ٕC���=*�r<�+�=���`�(	o��Em������v�Z@����`�y�v�I!:�J�k�V[Oo�ggs�����]� ����=Ĝ�&[�D�B� �-.���Х�iaJi��ڸ�X4A��:_Z����o�K�u=	�%=���_�a�kSmI�g\��3��c!!��g��������7��q����8t���ԙw��́"� w���#׵��3]	@�g�p��x�N��ܗ1�;�y\�.^�[�B3�;x>@��Pj���0� @�X��VD���
5��9�Ѓ�"o���5��D	8�6B�p������h���RY���5��/<��e8l�����<)r�'��%�N��qh��E�tl.�q���d<j�Ak��N���'�n,0�5�1K:�O��ϔ)!�pg`��AK;�������B�z�lhpО�;��1[�l�ku
��s&��?J��̣.���"b����\��h���c ��౳Y�4���-�A֎61 %kF1�S��H ļ��@�1�Z	��'�%�_�Z�w(������[C7�p|r�z��H 0l~QE\S@��XY<��=�9�q��:1�$�Psm>WY*�z    IDATG���{�
�^d������r�yzO�{��Eiq�rR���֐��|�;�i�|�V.�?��*[��n|����Y�~�lR�?~��n������~'���e݋��w�:s.g�[#IiW����X�d�c�M�����[���γ��	߇	��������������s;����_"G�4L-D��������4�a8��C��K�l)i�yY��i{q���/~�i��f�$�� 	��l^6*��hhp�t���'�$j��C�F��~i%��ka��9Oe$TZZT�֭�$�44rT�P��Q�]�s��X�m*�I�%�7��g���6�(�ሿ���2�f���ҸD�	����%�%,W�Y�þ��h ��<���`���@�7�Q�9�&s�0S�/�Pv|^�!���Hg:��k�tnSN;��3N���/a��J��(Mc�5nex�V!�Z���:��J�OL���)�-L�@N��E�*a�g�k�0�<� ��|��x�=QVX����9���;����K�ٝ��/W )c�أT��n���s;o�i��15&�EO���k�w���� �k�Hb^hlm�9+P�m���Z�}{��&d�����}�Cd��qt������I���
`�|�1�C(� uxӄ�Ȣ��8Wi��% `�'ϮD��;A�NDY+�4cA��&Y�L�"ekSIK��-�������L*8�Ѩ�bQ�A�4�ҋ���\BUVS���$ 4��?:���I�g�5M	%���<�E�i���!�_V�)O|���xM�9�N�_����GZqpȆ��e	�N}�j��p-�c�whiks�v�i~.�>p� g@��s�~���}$|e��j|�\%<�ȘB����y������,��T�M,L��BHպ��ح��ns�>�nO�k٪�7��:�t~�;�����ς����3N;�.����Q�`C�}�����?u3��6}�ǃ��Cl���I�C&�x	�㚢C(`�$#͗ʞPI4{x��_�E�ЬT$�x�����$-� �+��&���*G����Ǳ,T�?r�/�C�ݠ�dxg /��4�wBy):������f���{�]J���%i��1"��R
�$�%4e��/1� P�ঐI�ב��8�l�(M_օ�Be1�>��/IIF�3��
VF-���-?�,>�S����:V	d�{�Æ�/�u��3���.��?�iT��tu��=�(e��^Ƶ�oPl1奧YcJ�"�������z�2��;���D��ڿ�Jnd�xF��`~(��7_dS&wXGG��9���#�sK���
;�#m��l��P��>���ZWW�_��i2����3���|�Ս��X�l�]w�ٮ��Z�2u���d����<�+[�n��n���f���vԱ�ٌ�;��S���;�9~�T$��� �f�V �y������W�8�BZ��IҒ�*s\tE@�pB5�fA�*U�J2c��3�8�s��� @������Y���L[�c��Q�%pR2�l~� 'c��R�8�oi�G /�� ����ǪSct	'#�~��$��;q�S�=��+��se��)*��ay����D�`n%�@�DH3�Ж�Tm Y�(i��ro��i0���ޑ�QLX�N�̏��1�'��e%�]Y7D����;�_���w���e�"o�@�&��Y��).^�eoi�GQl��0��'ƛ�ZI�i)����m?s^=�Y��~���z����8�;�'�:�̳�^�T���h7��U_͒$'t�������{��6��-�gLJ����O�޽��=��\[�����`��q�-����U�l�̽���Z5	 �� ��(��g_�j�0�p�X �����E"ڠ�O(��Y��}Y4lp@P�,N4o>�"�cC
X ��h+���V	�(-�c�X��!�@)^�s���@ı,r��x>�%@����#��Cyj���A��{S�Ǽ6�(t# L?��H(�
!� 楱`��L���C��Q�r�ATcƘ2�*Ɔ�e�'�n�B���I�$�D�����q��K�zi�+	�f���X!��K�j���lHn+�J~����4��������ʅmʂc~�����Ip��!�G`̭, �7�Ǿ�={�����Z�E_�'�>�}A&Mj�� ���i��������v�gy�����q���zH�VͿ�̞3�������?�&ɤ�ɮ�Ϙ���������]w�e��l��EV(�ͧh�ۇU�cU[�v��=/��4��6��j�ڋ8r�E�_�$���~^r>k���=�� �?]����\� �hҮ�[� ���D�R!�A�@6 �6�|/��84��4{�� dXPb
��9;ƞ"� ^X�S[�����pGp�Mw�N^7��s�cm>�͙c�X ��+~zG�LƵDQ-�=��8�ZB�p��5�ye�r�1��!�$A]��;z�.���X��C�^� -
e��7�x��h��2#5b�t�Kb��\�ԓײ����y]�J�p]E�q���z��}]?��5�=뚦8L���/� ��Ų+�m����@����xɋVA�kZ�RM��E+��l��e���o����ו�{�C�6#�3ʺ�`���ȴ���OHh�]��?�{�*%�f*������t�1V.��E���\�i[���V�\g�b�.[gx�;rj������,�йP�3�I�������<�T�qj����7�KCf1�)�bt R� �~�3A4n�h@y@����;�	���U5ZK+���}i��>���3��{��#\�c�5[���ϳk�а��F�g\����b��������v���:4�l�XQ� �;Vt����M��jn��-?Ϡ"p��^ ��h�oE���s�K��N�g�o�%̽�L��M{�S+o �y_��~1t�
�y�.`d�# ���
�'%��[ ���Qx��|w,����σ:XÊ��3����}���`�ux��3ԟ�_��m�ݶ�i�;�g���"����\���y��*�zM���>��K.u*k��.o�l��Zص&����	M�t���\w>��F�?���g�W�{nx7K�.�g?���䓏�je�V�Zl�{�C͕T��u�ڲ�]68d�t���+��pL�����ᣄ���S� `Cv�a.���tg�Lhmti��4mD	iʘ� ��� 0c� ���f( �}�'��Nc��A��u�h��f)��}�B��0���1B0�q��b�Z�}b�I��-� ���(ʉ����k�D�W@�� ��;B� ߈�r�s)�|��=� c0�Z<'Y���.��� o���%�'�P�=��C���R�����o&b������{���w��?��2����p4�{��c�QV���>�яگ~����e�w� hտ�˿�� ��1��S��<�����;�C��Y�O�y����\���6�_�g�Y`����.��N�����������������hNa�U�o��Wv�y7{�{n�L�b^|�~�����c�R�׺V/����\��n]�-_F��6{a�:;�����x�ob6%�ڕYy�%�x/� �x�|h����O~�V��E�H!~ ���E�p=��j�9*��DE�<p��@y��@Bh�@(��P:�g@sAh���Z�|T����#@u�<��=��=TE��Z���O�TV�h8����|g��;D��S���`��F�W�NƇ�� Tm3QE�0WC>��������o�9繘/���،3�@x0�Xq�~�G�Y�ԍ����q/jN�Ys��P��=h��p4��p�ui��ǅ�t̖Y7�s��Ϙ����v�[|%���͚&G��o�����H��8����+���ڡ�c3fN�^���2�A2W�����-�r�Ŗ/�[�P��|쟼�iw�:���sYT�4��̪��c��/t���4�Jp2�������h��>km�ط�u�w�V.���e,�_k�����Z�Ζ.]iUk��K{m���eeX��,�h���7|SJ�C{@+���˜&��i�h�z���XXrk�� /�f� ^�L�C!�h���"U��o	�)�����������[|��Y[��u#�5��ⵡ"���~���M,���c��������\Cxa�J���-��y@H�G9n���x��k��V��Q���S�;j�uy�)kQ�g�y�x��!�'�h8͕H)&��-���	��	������ܷQ��%�K�"?��k���~�aW�k��C�A����(���J�͟�_��9{����C���۴�s���P��R��E֞|b�����_���d{׻�<��*��>�9[�d��q	>���c���ZҤI��w]o;n����`?���e��T���k=�~��,؋/,��]�mmw��?�-^	&$��~%K}�c��s�=�Ԣ��E�H��;��/[��ə�8�F_�`��I���|��L ���EI�i��t9ͅk�q	�Pf�d���Ikk-bHQ@�6����; �u��I�S<~[Z��{���=�??�S�9+UVL|��P����!h%��c(���z�}���a1��b���Z�2����\>S�#Ń��`�<��(0h���j�!�>t���H'	������׃�蟗r�M���;͹|=��1�>ڵ|.�h$���ކ��j I¥�3��V*�����ȦOk3��k�J�z�j �,�j�y�X_�Vuu��g̶SO=��i
eOo�֓���������[�\?^�tG~)C��?�Y�/�]�ٙg�n��>�z{�Zo�:[�f��^�Ԋ��X�
�P�����ޛ��]����Yg&$$B"�B�w"�Z��IP����ź�o�׶�����V\��KMX���(UPA@�%����6g2�Y��{?��̓Üs&���f�����[�����7R��n��$���]^���Z��c�5�h��[5�Ź�lX�9G�K(��}�r6i�*�`S�v�J<��^��xnv�h�C��܏�b�'�h��{	E#I��<�T��V��'����u	%�8�ǻ�X�����L� 
�8������	�J��w	͋�8H���w��%�]�KBw北�:�����d%j�c'&�AQ;ʚ�w�}4ǔ�@��Dsƻy"�~Z��0���N���(��yz���������/E-V�� ���Z��S�#ʕ��E֘�%]P	,ٺ�)۸i��ض�JղM��[-�����lp�j+�Zk[���eo}�͞}�U��~�;����l�#s�h�,��_���
��w4�} 6p�Cgۻ��v;䐩V���y���l��uT7������������C��N{�2����>�X�;�0��+�ʿ�Z��7����/���f��6��s�Øwf#+kT$�H��"�A��7����'ϣ�mi�Z�z�84��^�v���6)!$s_����eE+�~��������VA���&ca0�H��#�� ��3h���w���u�ݩԂ�c�'��X�`.8^�ɵu��+s�υ�������<��k=h����]�G�:��?~�;��W ��E3����������G��k\Q�����̄�rX6@�Y�YG�j+W-��+�yC�O2)UISV���u�y��c����`9���o�b�Q���V#�Ϝ>��ŋ_�8G��5�|��Px[3��dj1�ɋ^h/y�mBg���)[�z���w���k���-�-��ڬٳ�����{�M�p���¡B�P�MY}6�e����͆)Φ*��/�C�A�C+��6��ٷN�H�i%[`  ��x�7�V��.��K��I˽����J�����o��d���w���v�W�X�I8�z
���9�o��OE�$�~�Lڲ� e������" �oqss@�#�j�K�wZZ�Z?z�V��-�+Y\�x�Ю��s��Oi���9�_,9^����Z��U�,z�}4�d$���9w�(Ǘʡ�&3��L:G]����Ю&�p+�?������}Bg��c�s#��[��=��mdN����E]d^�r�V�^����,�e˖z1��g�9�y����̎:�y�7���w����Р�}=�}���;7_w�������P���f�/P�=U~�$���KmE���P�3��߱���cƌ�>�^�;���l����YX�~��}CSo?�'�E����rE��B=y>ORK���QYh�W���?���;�/?@��wh�X�y�X��CDE�rs��CWI��i��(��	�h�����|_�?�'n�g��Ϙ��V�Vi쌯Jr<mc%����s��BSS�Ɖ{ro���+��9
�9��^s�8�.�*	X渝e"�wAc幜���I�B�B*��y��Z	�X IK�����Z�\��|βD�O,������pP�J-��0�����)۷\Jh�&�ߘD��.<�T��h<��ݗ_� ؃zn�(� �v�*�%�O�l��vt۔��G`��#��b`����Z5�wt�����?�����B���'��?0�����.���)��w�PŇ�r����7�ѝb+4�����+&tǎmo��lHi�L:M+�� 
 ��[��V�U�`3�~������4�j���b�1�<<?��;�#ԏ���R���� Y���Ȋ xV��h�h� ���(�#\ �����w��g�TbB��8+�������e#K�f���bR�f=��k��}��)u\�1㠕ƈ�!��3��zH*zǆg-	LCƖ�b.9��C(sՐ��J��J� Z�"Ɓ
�D;�7��:4s��o~SO|��P���t�Ӻb�.������{�΂mZ��K��ё��M�b|�?�Z(��1ɦΘi���\���~���m��-�t�I�3����+h��+%G!��Zan�3{�t��"����c��;|/֟<�Q>x���e��X6�	�lGֺ:����R(��u&o�����?��;�Q<;:r������>c��nY��+��ߦ�c�[� kq�c�R����?����d�׿*&�����ʖ,y�^�%v��G|�]w��ݐؼ��ԅ��
��G�v�-A&�q��N���zQ�@�I ��ffa�0
��w�$#�k��.@Ģ&I�Qug ! _�HBR�H��
�8��1�t��3�q��V4Ҿ�}ėJ����:V�q�Xm���i�����T�&����g�4�'Y��	�)T�XT�[IZd�2~܏yc���/��a^G�S�Z;�Gt� n�e/{Y�i$��G�+k��^��C����%!�(%��sϱri��{�~�*���\&� �
��ZMp=��'b��Cմ�>�X�5k���6l�b_��{l�A覰,����#�u�%M���.�>s'kPY��Ε��P�s���<���ʎ:�9^I�=�N�c)�LV���ݕ�L6������ZP?��߮�;#m�IS�~�-�|���>@cp���*Ւ�\+S|q���I���|�	�I� 2|���x�� ��-FE ({Pe��w���� x��&͓{ΊL@!	Iڦ�F5o��`I ڪ������Pb�Ҍ��І%(��c�S<����Yisc��|��u��[���-򪬲H�)�ڌ��=O5c�Y+l|��f�'ƛ����an��5�B�C �@�ɪD�o���܊���=@���*�����P������������[b�u��V�Zi�6oXo}=֑!>�b�r�i4M;r����J[-3ѦϚm��j�j�
�}��k��ǟx�)��4���E	�� ֘񮪃$�]>1/���7�@F@��ɜ����#�������p-p�`��g�Ppq�[\�#O��m�f�*W��w�C�W(��UK���������B���>���F��
�;�x�5��    IDAT�B�g5YV_�R�/���2�/�i(����O�����^;Nk @$������rN㚊��Bi��(0�f/�Ţ�z"��De�*_E�x+��H�q�𾀓|	��POT�~W�6ׁ���2�5`�;C���{_���~�O�u%�>��@	2_rFs,Z�֔@a$��Ɗ��'|�o*�J��7��]&�c����r�s����]-�s��'�Q�xY	����?���=�[�@�M�r���w����趘���Q� �TyЬ<d�V���7[�Be��[��'/��CCUO�*��Us��9G۔��:�wz�_�p�=�d���!l2��.��b�Xrq`�LD�%�}�}�K_r˝r�u�]�E�"u�1��͘8U4y���o���PV^�*�?)��P�A�w�'���#��6�g���)�����=>��t�~ܙ��ģ+ X,�P��j�] ��OX��~��C��Omj 0a�Ӳ��f&���}��"o��3�i�5�U��X%�(�H}b�q�Qy5�V	e���`��,P����Uw82.� ϳbEȼ�;@�s�O}h?5$G� �|��/�k�\�Uc)*l_9|���i�K��&驿��#��
��8w4:�� p��\��^�U~�VI`Mh#�S���3�|�u&ڌ�#a�Ԏ�Q�'ϫPN �P2@|�ִ4����J�h�D��+���s���{,���Ƶ���c�ufҞ�J���~���8 תVM�l03��3�&M>���i�6��_���VZ'J]RZ=r�֚���|<ק?�i{��<�| ;�r.�k��}�<� d�3�Y
R�<d�X��4�D�|N�"~��}),�5�ã|�7B����Y	h���}*�g̼�L�j	��M��W/_$9,���31 VtO�P ���*�aP����������y�Q�i7oݭ�U��I!ڠ]��$L%TR �������� ����DkDp����y>��B&�@����;4Gq�,`��g��:��Q)��V�R܋��Se��K�_���g�]c��͏S#�q
%LT*�;|(�h�|���YT[�8�����P�*��5���fYc�J�MF�h�N\i���M��%��=�X��
�][%z�K�0N�Ԁm��rV�5�V��-����Ւ�,� ����TΪ�iv��ϵ��DK島e�v��k׻�c4�����?�'i1�j���O~�֬Zm���7����~ʂSߟ��1�Þ}}�k��D]ʊE�ↆBX1��I2����#���Jz�|�O�V�̘9��o���_k<�}����,*t.Q�'��	��K8�Ɨ�$c^�b�[ȥ�l�i��f��|i�, �8\����1�i���f�������s��sU�+�CX��N���1����E�v. �'@��@·
R�H��X�*7�3 ,q���� � (Y ��u�w���x
��DК��G ǽEY�V�C�Z�[\9U?U��Z(���������{	��h-1?qKF��|2��sJpKH�* �IDOi}J�ig9�{Qh��yN���i'�`��+C�~��c^�����ͤ�����A���?q�A���i�7m�k���=��S�'YJ�kY	�4Z͟{K@�;DΡ�S���N�(��0'�7��/��/�-Z�w�Y�A�Y򱐕BJ�N��)�(7R�5�T
ڧ���ߊ���-�I��a�g@��ed��ؑ�zh�f�6rp'�����l
�pπ�J5��]K�KE�p��.�f1�%\����z��,�&��k�+-��%
�N�)�x�[	1Q^zY>\[��! >��w�j�tہ��~��k��ߧ6.�)G�@V`�؈;����A|/ �z�
�JK���{�ΕI!�����R�RxX#G=S]�%]��.�x}����x.5�܃:Bg�q�k��r�i������W�N��.Tm�6�τ����߶�`_������K�ӹ �{��+�_�_
��]�� �1g�ׯH;|Z̟�nY�Z�4��A��9m���8vi���@5,�)Cs�j�[p�8O ��	bT �2����F@j�6��9)��'<���:�Mh	���L;�ԤM	|���:|/� ˃��9��:Ց��Ε�(^�Rڹ�M��Oi���j {����3~�����������v�Y����x��4F��"S~[e
�X��Kc+kP�1fXr
�%̹����@V�"��%4W$F����<�-��;�z� %��8�T�Ҁ��l��ֻs�u��CA=�\����;X��G?�&O9�JՊ;|���km��-MYD����h�I�/TJ{Y�1Zl5s��B�+|r��}:L�p�D��ĉ��aǡ�M`(��aއԑ��8���n�&�H�x�w��'�$uК[���~
��EݼM4yi�,8w6���ht6�6��G��1�h�I𝀸t]I,��2��'�]i�a�,:������������g�<���qכ���5��[�RG��(�4 |���d��=�y���%KB�p�rbK�yD`-p ŵ]�I��@?^��;vr{�H��²���Gkݶy�-�ԚC����gX�<d��۰v����p���X�])��C=�ռ~��6��Éذ-�wؿ��ڒ'���	�] ğ�̓�	u�g��-8hC�����+�H{/�S���Byaܓ(�B:���q*������<��7[��}�å��,�$��'��A�%����Z$o0�[�n�|E���<S�x,xb ��'��Sa�X[�5���y��Z��b�ǀ��γ
D���Lև�_����k�1xb�ƛA�I ��0�y&(�_�>�<�1��V�A�q���X�J+�/f5�r
�u� S�R $���� ֕����K1�wAP�+���V������4�����M|�YgZqh����n�`�};]3�=��}�zy�9N��6���6}�LO��oL:\�f�lϱd�j���)�Z�{SV����֘�Ա%1]Sub`!���+K�-�,�$A��l�q�g�U9a�8�����3�N9�6s��I-Z�9ߛ$X���]i��9�L��� TG(:=�|/�1��c��5�H��4�F��X�-Pӂ�~Ah��&-�V`�0��5��Jck|T\_QJ������#M<�}bMZ=~e�s�6z��^��K�Z!v;�hT$�֐Rc��<�^��敟��@9��)jH�C|s���ח/G�+%{:��x���8�=�7e��;�s�\����?�{$��p~���/�L;�&M����t&�͈z�	�{y�x]�oQd�?�B!�!<�)T�$V�4�u�<���%�v2I�"ǖ� �#k���Z�|vu�����g�w���74����h�6�_s3j��OU��i�!Ty��uV��qG��	-�����v�g?,��Q �w�7���s��cmN�/KC�F ��,J 8�2����%bm/�$F2y�1�Ij��D;�D���p��]}-#Y-<���B����I���S��4�=�UP�B0�!k[m	�T�:귣���+��w ��� �t,e/���;�Xo�7$r��wYd�����w�q�\�g�6�Xu�O�g��?����Li7V#}����֑�oϚ/-�U=т��"�R����rŲ��l��e;�Dh��YB��aa7)B̑�]މ1�
e�Uԑs�N�_�ּ�0��lG�[n$l�P��;r!����CuR���X.��a��V~��X�o]�!h�>95����7&o޼s��Shf�8�7*�*��v����,&Q�>ͦ�?����c���wo�Q/�&-J=�x��ħs��?QA�P�֢��(��ck MK�]G�[�}�����^���zҤ�;O�2�}M���K�$�s��]*$��*5�ԛ���n��;���@����_Q�� B���o�ݣ|h������������A�A��AV)돜2K�l~��_y�!�{��_�E�PD��d%��q�����T����	��Z�W��Z�����%�fRV���9��V�f%�}���Ý�MI�0GP�t�J���aI瘮��m��J��+E,Vd�/�r(Um�DҜs�Qv�s����&L���*p�|�
[�jm��9���wtUUh�ߦ�[:������zgʪ��o���E6��s|B���r专�R�y�Q������M�;�(F�W6�w�i_|��� n��f/�,���B���&Y
�}L�H;�ƌ���v�V��"���.��G��o�L�*$H%��]�P7)������J���4�%#� Bat�g"ڧ�;P�3�$��'���_���l"Q���44�v ��ݾ��o{���.��rX�4���_^_G�]w���34a\��^�'����?�����ČG����g����̥qݱ��B���̕j=i����[BC~�u͘q�W��;�8�y�t�|����{����k��ҥ���w��a����;���g��i�r�j�Z�>c�{oY����u����-4������P�L>lj�ܜԩ�_-��n�L�^��/8ߦL�T�����n%�~�͆d-Kel��^��^���1@S�����\k#&�l?��O�/x�oR����ы�Q�)iӇv�&;�H&c�s������Lp��( P.1>�`�w��OL�	���X3���{�񓟺P�v)�E�.�&1�M{!5���a*���E�A} (����J���??h�q�>�nD%��CH�������3n��F�S�r l`U��J(X	���Z�b$���7�#X�?J�����|��|�7����b]q��y���BG�&�\l5ǁ���������e>��H�ճ�/^�:[��'ͣ�"X�V,��Cfx��'�Xj�/�D�\G�	�'	�#����V��Y|�^B6oC��v޼��k_{�M��e�tնm�l+V,�%�?b��l�,����c'�x�}�s���ȍ�SA������/4 �۩�����}����Q��+��K�,�ו���
HY,&z�"@�8P'�W�d%����v�F�l^�W� �>��j�/0�3���[ns�U��w,�Z@���)��wн���)�����[֯��3|G#X��<�ǀ?7E�����}>��	�#�i�A) ���0(�} o�h�����6�( (%� ��J,�������}3YN#�5�w���Oh�.���_�}�dK9����U=|QT�O�-t>���4����VX/eֻ�y��m[69��!3���͵l.o��Xg�{j�*/'�z��?�h���j.��_��?
=�����3h,@*xN��f����J�1}�UJ}�}�f{����򧞰����iV�x��!���?��<{� 6����
C��_�����|�+�G#$=�]W\�<-ş����E��i�b�̵`�7�E�l�V�C�����_��o%)�`���i��Q�	�"�~l�[n���q�u�G���FZjD�#m�����?vFslɆX����G��\�5�wu.c�Ӵ@F ��W�(� ������d^o��G�G�W�.���_K�g���w�!����*Ҁ?��I�0N����D���O+��{���"�u��g�������÷���>�N�G9 ��Cq���g��H^c=#�����g}#�K�?�7�\�Ry�{�a��{�9�Dp��6�?ds�e�}�͞��x�G1��n��P
����9���M�r�8��T_�k���۲��-y�!{��-��zQ|fY�e�lgϠ���q'�j��z8ߗ��e�p��{�s����I�OU@z���	ƥ�H״-�F����"t ��5�q 	��f�NL-5�rů��*���B�i� ɢ�;��{�}�����K.�gD�yN��IS�ZV�,�}�9`�{�+���gV�Z�w~��c���9����p��O'1�D��{����h����5�s��� a��������s�T��5��;�cF��so9|��C���D(?�e8yk�>��p)#�1�ozӛ\������[xXq`��z%k���\���sө�elȖ.{̖=������i塢w��첁����؉'�f��y�z�,�,��f_3���4�����k�N�6Bg>o���]��c��T�h����6uY{�l��^��R�����l��-60h�ik�����y�?&�g?��kq��1� L�/~��&4ϸ�7���dS+$NL� ��9�|�T����88���� ��^롃q$�H�B�����1@?|4e�#�U�(���h	!m��8��m���?��'��GGçp��>����zVǩ���G5�YNz�/s����8��P GB�n lE}iޕ��#Q5�&c�H2��(tX�c��q�OE�R#�۽d��u�gl'5��u��CNH ~rB-L�o��?����������h*X�>�j��p�c@����f������8�k+�z��%��ښU+Bu�rj>7�֮�d�}CV���-o}�<m�<���d?���u!+ 큫����U\�3�����:<�䆯~���O�\�+��_dCfҝ6�_�IJن�v��'{�*@ʅ	_�0A6����*@,�0A�C[ToV6&�P�D���׼�����PWg�h��.\���V[�xbU��u�<1M�E��_�!��K������V���p�bR�$9���x'�h�h���sEg���
e�. �xʿ��}���.��r�_EH�Sf�d�i����u���h����^q�hȝ�P4}r}��a�vCͲu� ��m�\��5s��w|0�l�ga�`�C��/ Jڗ��%�A�p~����ۻ�CgL�I�'چuk�FQ�u��r�f+W��J5c��vۙg�k�{����k�-]��n���m�������T�s��q��?�c��Q�~۸a����;l޼S,�.���Ox�_b�k����m��V�u����l�	��#���&���|����	11�x �-�_����:�JQ�Y� �Z���(K0Q4\0@����<M�@��qBSi`������Y�ȝ�q���]}/��������D�ƅ�u��1�{�IJ������<��T�����d�ǚ�(A���c?.���j�����Bz1�-KNV�֔�Y���؃�����E����$vՂ �4�g�c���aܘ+�p� ��ĺO|���u��,p��"�/���l�#��_��N9�h�1�[�أ60��� |��@��u�u{�uvM�_�q�wM�����ƛlŊUu�����p��3�������o���>Գ�毥v�s�t �Z�V�z�~������n�T�֭_i�}=I�D��-ڪ�i�m�/�`'�r���M6�wh�C>�4z�^ >��?�&'�mTB�LR0L��E�z���d����q8����Z��Z����+�tx>�Ef2���P�lFۇ�G�W)�v`?ҳ ��>�J5ǆ��y���P|�`��)���� 4�틠m)�E�)	7Y��W��9�k�B��6�Iܞ����z�XP�^��i�~��n��KV��^�*[�x��k�c_@���o�i�J��;o���8�>x��Z�<�zz�0 e�=���Ga�v�����~β�N����o�b�r�	Qy}Y����?_ڬCg�'?�1+�,m%��o�h���ݶy�:��� S-c=�A[�j���Y۸��iej��ѫ�O�����L� q��lp���7;��������ϙ��)�ub�w��A|���3�n�k9RZb+��H�w,_zH1�#l�/>#�p|�a��d
)������s�|�|4�ǳ���c�Ɖ^��k�ɇ}�u@���k�|��������5����N��`lEi�]�u�N��'�G��6y�Tۺ�ە�U+V���	l��������w����1k������i�{���}�v�
+��i�N�mg^��v��m��m��ګ_�jN4    IDAT�z��=����N����F��w^�.����)ޜ�"
ɹ���8��e[���L��4g�� J:�xB�	x���?BVj>��Ku�#�>�x�!�G�/*N91����N���������=�C�8�g�b�;��{�#f�Y�kV�p �8���oK�\a����M������ezh���k��j�=����G��V��τN;h��v��U�Cֳc�mߺ��wo�Ri����%ˤ��/tÆͶb�FK�&�;�����~��1�h�$[a
����O,�,e������׻U��H��J�#�x\��}�
b���8rM� I��~��	��磈'ێ�!
��V|SK��n�������ڱ�{L����C�N��X���O�Mq�*CQX(~�;{�R����l˦��ݽ������}#,c]�{G�=��%ֳ��.���6k�l�T�v�O~j?��-����)��%cx�:|���QU�t-ms�εw�������[��=��a+�l�L�f���@����c�©6�9�8@������$ƟJ���DD�"5֮_��f��0��deӡ��H����?�m=~�31�p��V�+ �Xxj�  T(Q�s׭�����G�3!���c�1�X��V�]��ʏ}���O}ʁ���\'J��N�qQ���8�@	�_�q�h�V-�e˞t-ʇ��\�_���`�N:�t�{�)��uX���]��=� \j% �8�VU=�VO6D�,���)S�S����V��k�����k˗=�WS�5a��z�iv�9���鳼�@Ov%�J���D�/Z	�-���� ��N�V����J-s���7�5d�9�q��X�l�+�EV �1�OTq(t��1M�HłA����9���,h��<�x �XޓwW4�"|ؓ���<��x�c#G0>u{� }@��˟gR4?��=^t��T��Ѐ=��v����+�[�J^HH�<a��v�ة���5���<��gw�ү����s`W�lQ�_]��JE��5�bG�������Yg�n�Ҡ�je*؎�[��[��'|�t�T�e;�X���y�ų�0�lU�'��/�ω'���]D�ȩ�yh0,.�>o�1���h�fe�h���]���3kmK����=���TB��b�e��T�#�u���Z!����eK��iU��ݳ����Z�]�I8�	�&��g�P��������,E��	=����ՙ��ނu��ڵ���c��>X3gf�"��t�._f����~ *��Ƚ�g��o��Uw���(�J}��|_����/8ߛ,PB�hRJ�ԩVC��޾�����=U�/����W_�@�ǂ���+}�X����_yHQ
,���ĉ.��9�� �������0�S�-�]�z�gvS���P�b�W�H��0�U-�N۱�k�$B�<���z��р|�cT�	P�ު�p����+��Q��`�<��Hй��P�^������_w�[t,+��~����o�B��G}ܾ���Y���^5�\�~?�����
݅KGN�ҿ1��o�P+�F�&L�I}��W;mCyg>��eaB�l޼ս�j������1hj�v���A$;�ݮ����¦�|���f�����u��E/��pdƺ)Z� r�YH�m���RI�K~��a3C�ocl��Iy�V4��s�єw`̈��Z�ot�kG��hL�	5T�ߎ���l�ќo*9��7~/@�3�UnC�[��O�c��*˺1���F�&�4@�������Y:������<P"�s��@V*�uMԏ*�����^U�U����Ο��:"��G��t\��ڱ`b/S��w��l ��_Ia��vK�N^ټ���!�ε��&{73U�,�"���3"���==Ng��O�������3�?�{U�er�w ��9�|SQv�֊ ��kA�����z�^p�c��G�'�hB=�N \i��$���MD��JU�z�J�1h?�z���ΧV�C���0S%yQ�ᐩ�F��5K�P��| ��H���I-s6�j��o�AJ9��y�X9�v���PVl�Vr�	���v�h�}�{�kK�� 9�5*�9(*I���<�ϕ �2ʄf?�0�}�o��"⪣�KZ�?� ��GQ�\����C�k:�=y�s	�x���8Fu���
#�{���zdN��\=�����I'�uE��1.���}^��н3��gýR�`!��F�w;����߬\����!�������`;�Yw8�� R�l*d䖂êqQ�����'���� e`)���O~�K1P��k0���Ь�Z����uY������/��K<;��z���$�8r��w�'�2��1�uI��nu�������f;��X*!R��#�*!�ZD��9����ƒ{��۝��R�S_'I��:�\IJøގk�{��%PdQ�Y���M}�����E7V�˳���R*����7�(��8�X���r�����%y�w�q��ؒ�] ��v��|�a�8�9����&�KR���_ʹ`���Ă�n��(���;��2�j(՜��10��hh�����©q�aځ%1��W:�����& ,��iQG�k�$��(
M��.����n�4��q-� ����S�3Lnh�^L� %�<cA�CM��%%,Ne3rV	��B*Z�#-���H���i�����4��y󭷸�[%k%�)M��c���;���Jƀ��&�*�;�I<��6�~�r�&�����+n��F��I��=�w�y� �`Zq���)�����gkw�-��땠Z�$9�S���Ny �͟�J��/>88�'�h�=�H߫���Uq,悬b�Q��P'~R������:��4*�uKh'-i�T�d/�I���z�p��`�9t���c����[�a����:|��)�<�n�jA�G�
�t��b4�J�ĭ�r�w&NG/��D�o��w�Q�4p�	��4B)8~B�`�?=}��\RW��O���P�v��1�ƢVm�F�_�E
��@ʂ�7l,0�	��ӤƋ�Ն�����8|���t�Q?5~D[�n���$� -���/�_�\��o�y�V�֧�㿧�6�S\��)�d,��1��3>�C��D���1�ז����+�Hc0�wP䞔Q<�p#t>�񏏘������j�!���ZA$��t�M'�%����.��{/&��?��S4vj��9�ƨ~��0��̹j%r �p��TI���F팉Ŝ��o,s���v�]�a3�q��D#�����y�E���c�G�̹^��_���GE� mC�&	o��%���9|o��mN��;�GμUO�}|���ռ�, 61�<
�y�ERu�&}�1	�?Pn�~ 5�6�Nh !�^c���7���X0�bJ�k��%81VXI��sٝ���c��Z��<vXJ��6�ؖ���5��s-���}ޑ�Wt��>��{����M=���s	����#���[*%��L><Y�h�`����j�P�8(��c�lοE��k����HӚ��L#�j��PfA� �Cㅴεهs�h8��f���3�T�.�A6h�Ī��x�K_��_o��ݛ|���}ڙ�.���K(�H��_�����YG��ӈ7'�}�[�����Z�%�j����p��&��r��`����(��7�_�`ų���ʺֆ\H��Y��]Ig�� σ��:�hr�]�!a˽dep�7��u�[k�v�DϠL�՜�=���/���Z�7���/ņ[�ַ�o�(�MhY�g\v��۽����u|/�E ��Ou���]4
3)ij(q����^�B8y��� �]���B�'��F�g}�}�$�V��6(��������J9h"����kv.�E�*b3O� � Z���j*���U��lp	��h���z�����k�'�3s}@�{�N��h
�-	gv�Ӝ��J�½�������v��L�,��rSI��	-z�	��d�k�	,�m�=�>����
��y�K-�f��ˢE�p����ޚcͫ�|���3��:�_|�cu
E���<�p}���{�ܘ�z�K]KN/�����|
l5�;�m�Gćs��#k(���k� 5�w���5ͳ�}�� �@D�����}���,��U��4r����a�N�c�}��Ĺl	�f���]g�aV��%���ש� Z�j�qԹ,�봇4�X��$���ڔ�`k3K[��N	��G�^���":���7��ɤsP;�m�X̭>��X>ZԊr�i�+C�N��X�m�ϭ1ֳ�����Ƈ�cݐ�G�a�k���W�q>
oe^Y7$���_ �O�'��ց�ќ���F{���H�VS:᮫� �(d�1�K���G���{�ð��OJ�H�5d�"n߮��j�����5(�_ᥚ{Y$z.�����)+V�\:��[�:��0aP�p��q�R���bZi����Z�UfN���ŋ��5�I��z\��n8\(�Z�f3!<m?PA�
�d�<p1o�9d�2�����[2��P|���^��/ ���r���AlA��'`�l�*D��e��iNc`޳��c�T>��9d:k|��~��e����{�U�k:�~K�.��2������C���x:LUX��|��zA�v�/���g�9����E��e#ϥ������+�|߯��u�^X�-���W8�j!J��s�,)*��%�yX#t��3d�Ha�<�Zk�fَP�'��Tj�vM?X��/���l` 亠t��������fQ'�_�iH��gsA{��ET*A���	�삏/�dtuM���m�G�X��Y��5�"r$)����`���18�`k�O����o�������c˪����6
���v�?��ey0/ZC�B(���ؕ@˩����X��<�@D��Ɖ碥���|����xʊ�T8��=��كs�!��}+�_o-�.�ZPb�v�':_�[��["�CG������mw���g�a�C�JV�r�k�o�	C·"ɔ�r�c���OP:�Y�Dw��f�h,;�����eѢ�5��[��2�vH�pS*���<ҙH��#����zz��9��*k��2��7W�?G����i�P���c#$X���A9�c�kԲ��Z��z��3vJL_qSi����3n� V�\4�.n�'�I{$��a��r���D	<	t�ݓ�.}�.�5XG_�����+ϱ>{੓���[N�Ш=|����,���-T I�5�kX�D�L	����eB*�sR��E+A�č�[�#�	в���i5t�#�PX~ �O�?�"��-ʸ��Q
�|H|?�2�}*�O�4�'�@`��P�	��3�-4��#�wIݓ�u���{����I�ä��j����+��+_��L�4w8IY�h�ī��� E P�����P�Z�5H����t�Ӥ{���6w;�2Vڧ�{����힯����^f�45�9"����ii)7ɉx��7�R`�M��m6o�E�p} �� W��}^J�gQ�I4j�l�r���+�%A�t��(����^���{��QC�lҫ@'as׸��e�r{�q�^lq��aD�o��*�u��-<�,�o�%�޵�M�4��e�E�S�vJ���B�ּ�1��=���g̜����{�N^0<�=�Č�8a�k�z��k�>}�o.����pg"���r�
���d3�������S$'}�{�sm�c�S)��G13�Ac�yGF�D��]�����H�c�v�>���>#	����{����Ώ��;�M���T�t~�����Tkgo�"�ⵡȣ|�^AR�	?Q(�$�Y���a,c[n�3��ц+f�|�.�G�A��E����vy8���o�����w� ��h5�/zE��
��=Ĺ�o�g��	����,a���7��N�����3��a0��7�a}�\,��_����w�s�K֟�w����s`g�.���B��f�?���W��Ͽ���/�x|_�I�>�>��p#�-]�G}ԋ�!��X��$/!����!d�&�DkPן��4|�\���`m�FN�QP�u����p�÷Q���tO�c�v�����������d�b�1�lf=�z�{��^=�}��6����@��8�����J���k�j?Q���U��N�8-����9RO��:���^��:�SW(v�c�˾dL��ȇ�ͬX���	����n���d_��?��{�'��"�:�'|ods6y�A�y�6�ݸy�w�A��r��B#���m���5c�R��l޼y6�E^�&��o�f�
Ϛ���O:�4;��6g���2����#���7��<>���C���?����?���Ԑ4 ����E�&QO K��'5�ݱƺ�������C�'-p_ܿ�5�PX+hb�����x�����$�v�s4��2�&`"��}�)?��=V�����}/�Cs�s2Vʒvn��|
�#<�2�I(u��'��4y�Y?��T�z[�:�X�`1P�ΡW�%랂����~�m�C��W�%σ0�3��/���z��1����_�Z;���B����mt��rQ�4�����$�;\��Kig��8��3���[�F�$��Ϝ9�.y��v�)'Y�4h=;�ۃ������>!D��P�{�̙��9�γO<�r���o��v�Oux�I%J���ϸ��`��ٞHu�M7�BQ8� B`o�v��@��g�T�)vp>s���TH�Q����k��ۃ*2{�;�a'�=ޣ[{{lӆ5V跮���xJ�V���� �P7%���s���I���ȭ�
�쩕��uBI �	��s+�K|=���uS�����\P����~����Q�KKz(����g�A4��fO<�����_ن���EG�;����K_�J;�i�����3�����X�Ԟ|Mn5%�I�����=2gh�^���eo~����X�V����Gy �Х,mIĠÎ�ݶs�l�}�)�����d|�_p+�L�^ij�	��B@K 9�@	"\G�9ƪ9�������h����}������ڶ?%�N��J�^�nmw��|���:f|x^�8�qکf����{mӺ56�W0��)�x�\y��@瓊VLuج������X:�a�6o��v�=��ɤRR'��w�e�)���UI/|+�X�m�v����*��d[�s���N���?�K��m��'l��mǎm�ˇ���ض�������/p�'yq����5o ;�������G����f�?!��\Ʈ��]v�	�[�<d��M��a=�M�a#NU���P�6o�j�r�zz����y�{��o��>�
�BCIJ�FS�o���1�X�,�}�����4�i\��7C=�=�Cy��}"��Ya9��Z����[��P�m^�����[6U�t��QT~<�<4)��>ڮ��N�YGk��l�|�mܴվr�W폏>�+�N8ޅ�nr�%j���|�9�9���|��������+}��"��p��|�	�ʨ8�g}=�m���l˖��}�V+���O~�P�f����[�k��v���d�Ϛ�>GJ�C5������1��/�����U���#f٧?�I+ؤ�v����K_�+�ؚ�O�P1�Ϥ����o�W���!�������h�+W�ts�E�v�$oȞ�/QB����x!��(7I�g� P̡j(5���������)��=j
:P$k�}�{��u��V+Z�<`�6���m�,[��UܑN�r�g5�\��8�	�TƊ�)v�Q�ڄ�S,��t���7ڣ�?|4%v�ǘ��2�����g�����'?���wB�����>g���o��(~D"  �t�l���;��C��	9[�f�����~����mɓ+��s�-}r���%�_��I�z��-[���4�.92��`Ⴏw
ok�1�s�e������%۶}������i�t�֮{���{��e�����    IDAT�b�o�������csO8���	��/���o�' Iߑ��kV{$�LH�\�7�����G��J�ߛw���G@�}��Lo�P}6Γ�3��Ph�r;��ӬZ�L�d[֯���sT���x!!���:���9G[��If�[�q�]�MN��5�p��c3�PO%g�X[�k��N�o��o��ˇc��K5�T"�pN�İ[���_���v�I���i�l��%68je��R���\j��D�)XG���G>�e�=�._���ڨh$��f̜��3���7�oo��cY�l�a��UW}�2���Y��������ϰt�h+V>i��`����m���f�&K�'ز�[�O�+�����p�0���D�Ш�Xl��p-8@��r ���`e	s��8���z����N�V�K�z����1���Ͼ`ݣ��š�rѶ�_i;�n�|�h��̥�g=�W�x�������?�c�z�6a�:�_����ǖZ&��������/'� ]�^�erxN�{��]����T��}��\�(�|���=���7?��O?ΦM;Ȟ\����RC�\IY���Ǘ��J��ne�Q���������W��ei�z��
0�q�o���P��c���|�*������n��[���e��N��i�2����W�uk�8�j�v;�Գ|1�0�pH�R"���p�͋�uHn�{��_zM� ��Xi	q�X7����f�����5(�u�����1߯��S-�\�߲v���������<�����pNJ����MʩSژ�+�.;�����I9�a�6�{�I�>{����w)ɐDټ�U��K/y}=�����Ɗ'�+�6��|���n�Gp�Z��~����I'e3���_,FLeϜ��Wm����M�ի��f���_J���E��v�?s���,^����1hޅdls��9�=퓵��{���Gl�d��J���l��2��l����D��Sy��9`�W������ۼ�^��=1�E�VOU�X�Q���5k��0��;��]w��G�@ H�h�1~�����2�u����kd��x&�M[�0k^e���f���_.Yy��6�[e��[-�*:���s�?r��-D�0\2m�s��	��t6���W��	���h5�8zF���ڹ��m��]ٓƯ��4���>X���Ϗ|�#^�{�f{�ޟ�ԩ6m�[�&��j�O����-yb��Kۺ��N9�l{�%o�l��Ճ[�n��>�4���E��,DԠA��Mo�y�βJy�V>��OD��MV*S�+0qZ���wز�k�З���>��?�~*�+�-�_ř ~������淿e+V�p�W�Iu}�Q$������ZV�B��~�8�$�U�V�+ئ묷��&�3��]��fB�$J?�Pޡ��Z13�fqdh&di���o�����%K<)ʅ_�#@�Q(�(�W�J�ñ?�[��Ź������bG�9m5��F���gj�fգֻs����PiЊ��z��T���A{b�S�}G�]~����G[�����.[t�b����w8���uj��L�,X�B��n,��90�9�ܳ��^�5��|�=����z�2��-���UB�g&�����)���'�EA��?��?{B��_u>N?�tC`Q@��G> I:J�V���D�rm�6>��`��M��@M���ζro��};mݺ5�ӽ���L(�P){�j)�����[��pJ�lαϵ�3�r�fk׬�k���_�[�t���bv�m��b��GV/����|x��.��"O�BK��Q��i��fW\q���u[G�h+�z���1��3��8M^x���6ڑGg��=զr�z������
�Й�f+���)��Ќ�'kNN �-o~��ܼi��rY{쑇��?�gO=�ܵ
�M�2ɘ�SO9�;�X�0�5��~����U�a��kQ��E/z�O>���'�}�l��yZr�&ܳrW�?���bT�=���-��sfϱt��e��n�s��8��R&�v�5ۤ�����̆�;x�t���ٯ}��v����Kg3^<n,���Rv�BV�s�ᇻ�O�{��6n��A������ܕ<W�pL)���~�I��mp�����>۰a��{P�3���Km�aG��I[:�����{��7%� ���?}��?? ��/X�`qw���f௸{�e�v�An��>���b�y�F۸q�k�8c �9�g۔��Z���Jռ�%}�"����,t9�X8,~QM��n�A	 -�����Q���C�G`�G@>	��؇h��K�������i���JRO�`;��7�{�dC� ��syotB��2Q.y,�P^Y �[��f/��#�K}�TЯ�kO��
@�Wƾ�J���[.���'٤�]6��ok֭��[6Y�@�G;utu�o����������sg��46l�d]��R�|���h�\CA&�:�d�⬁�g�,jF�Y���-W�w�������ކ��rI�Z�B�������� �-��1�ݻǘ3~�d�� �>�F8�N�T��x~��E���?OS~� ���b3�\����/��k륤�m��nr�q��#y@�=��I�1��:�����_o(٠�`a�D!,:)�X�0V8f����^!����S�W��6�Z�����Qb�4y�$��N=��<�v&v��8�H�K9�t���v�]��D-R�	��#mGf��'���\n��Vw��!��}����kk����
�=K���c���n��ִ�Ls]V��U-nըf.O�2��}��| ��<��$d�f|o��q�!��)��B�k���.�GA��=��c}c��@_g�	�N������>˻{�96i�D�˱��W�xwa�=��?�w�����������颜�E��¥M����E��rJ=`�Qga@�I'�d�6+D��.e�n�:{rٓ�uTke?��^����|���������Iǜ�$���/}�^�{�g�������Ox�F�9�:�Gh݇it�x6g>��TÊgv�(�\:X��%}�^a�����pކ���z�*�M��aһ���b�Ja�h�T椌QK�ݶ���H��[n���<x(�SԮe��1Ӟw�q�QC���ֺ����I��� ��Z2��g����i��l���-�wh�B�K,��*�)$ӏl���W�&Y�.���+�K�I}�At!�$�aʱxT/����Z�*?�7���l���z��T���(?�o�G���V�F:sU)��M��Ϯ�<�(����@��Thv��tٓ���t���l�T�Mq�q����.��K�ѽ���5�y�G��H>�},���>V�s�\.o�	���A�� 4h3h����i�jq����=P��Z:|ہԮK��z�g6U�V�d�0� h�w�����/�ܣ}p�7 �_i�m��6����ydA�:_�$��03�}g��3�v���iQw��=I�zvvҌCᇲ�d;�c��c͓�"q"���n~������s�]H ����[�s��J�(t����9��\�<��Q�~���Iڵ��8nMg��Ww�ۃ P���H����8�"N<k��W�pfL��������t�v+��N�'�^h�� ��&�|�6�I�Rr����gqxƐ���
�5{�Z� ���\(t_Ҍ�i�hw�4�H�HׂD�F8�QC&#�i�${�(Xh�p��?�� Q�8mt9��=��,�F�R`���H��I{�������ꫪY9�Te3N}%�qR��"����ZXm ��3�;�Y�A�|b*�N4�D(Ś����8b%^+í��÷��0�`�?���`j�T�H��r+�|>�A3ޟ���1���F��q���u�b�|��i�E���@0r�E�m$�4�a]�8Gxb�oT6C�]��� ���[
݅�5�Ȭ�al0����ݵ�P�C��&l܀lB�b��y� H�ูs��_����G� ��|����ځ7k'��c�s4�����"��H���6����|�p�5J���F4��Q	u��Fo��s.s&
A׌��Aɛ	��g���]@0))�b ` 2����
�9K~�z�9=����]�曗@������/З(��I�S�%
�5��`sW���� ܓ�I�fb	Z=�����@���v�q�Ջ�)��y���k��U[�8�!�����hB� ��ڰ�$4^��a��*��:̀?~�x�Ŗ � ����b���;��š�qmX����M.����7��4���f�Цiw��o�}sd��j�Q������
i�~�H#��$:�g?��Gy��G�^"�D�i�wը?잼a;���w���e/�g!_I��Hӗ��"�#����<)%Nt�~��H���zaTJ��y�4�yXL�7n��S)XJ�ЇW�SFN-�^EK�okĺ�?�,�?��<h)��g�����������w A�5�@2v�{�����o���/�0��X��'�ä�$d��7"rX�h�Тb��Do5�rI�m#!�nc����O�n�d~�k��'y�]v��#�S����6��V~g�5�׽��노诊3��)ϭ�h�Q	�=��9</�Bx
��1S?��K.q ��C�(nY<�֦�T�?�C���~�v�d����� �IɆ䨘�ј��\���`l�I�fi��.�b�^`� Ƣpȕ�В5m�����beLc������0eLe0�g��Ɋњt��,��c�. | �u���8�9o�[���mh�с�������<�MT&�DX�p�C�x���x�Bk�)�����8�+�h�l��*i�!��NDD&�z�}����uɌ���{�J���ҾΫ��"(ش*�G�Y1���ַz��O��]�W`�����2�5XK��r������}�c@V)���F��H0��#Ǣ4} ��������=w�W�����Dah/����� �m;��Ԧ������O��ݿ�m�C��<�( ͵�K��i`}�=��z���X��t`�f�i$�W)_	�0t)��`ķ���8��bǵs����G��kk��%��1	!�D��eq�~� �`���h	���e4�M8���&�o|�;��m5L��Ip�o��q��(�y��۳�c�����$+�ͩ�
�CV�Ýު��/j.Q�Ma�d�V8����g+A�O������$�(,Z
�9Gq墴(6ȹ|�(�z�?���τE�j�b��-�,}�CH'�a�/8�����]�v��X�$�R�4��ź��[5�J2�+��#h_+Z,�V1��E�P�%��1pBkС=�C�sW�u'n�^
�<��$�HB���{��>M�R���Q�X�������^�W,�i����6|aW*aMS-����r�4�7���A,�4��c�\s�5u��V-$�<�?��@S���Vϱ��٘�?�,�GqB�G�d��%4��[h�1u�9n��G�ٷ�v�����_����Ų t�	�(�9�:�/�_>Ɓ�~��փ�����pD����빗Ʈ�4���@K��%��"��=�&9!�z�g���0Q���[o[;	����FzW������*9���`Q��^ba*�w�Iiq�I��	��  ��
H�s�o8����U��g��[-�z�q�V^�_�G1!Lrp&��X,{�	���PC��s��`��g��!�h��ڀ7�i;N]����5r˼����'��x�R��OPS����$υ���UO9���M�vϾ���%�{wzI]4���6&sR.���&��8i�Gċ4�Gy�#4H�{����2̳��4ƌ=��C��/}���������;�0w6�p�����w(,E��x��~|��O���1�� bE��p8�'��P@x'~g=b!���3���|���e;�Ph���)�(;�	�q$�F�_L�2�ڇ��~��J��E�J�c�j�;�9�5�����go����6���˓!\�s"Z����!<�����۔t&Ҋ�r�'"FJ�PցZ>C�%Ky"FH� ���&�����L�R�Y4L;͢FHk�f�x�21�)���SO�%�i���������/: �>�E�
`����6I�wؗߏ�1���	E�0?�6m�wN�]xw
�Q�	�j ��Z][��\@IQG
���s����������w��T<�a�5G=V���U�6�d<��z?E��"��(�����d��iR���Md��L�X 9���=���Xʖnų�7�F�  �<Y�R��(Q��bv}�Iu�l�f�:��BL���'����o�g�e�j5/���nj|@��k.�vO��&-.��Ҩj� ɏ�3�K1�9&d�i;�?�6W� k�5��/X
C#BD=V�XQ)--J�G~i.֕�;@qJh���Q@��&����m���x��Jh|d%p<�+�z#��kd�����w�6w��	�JCܟ�'���?��d]�����|�󰁪0K�ħA�1Q��X�_@��KE1�5[�����+SV�q�s�����$�+P��8���z&t�_U69�DU�a�Y��,+1�z6����`A��C(���<�1Yj��O��u��'�d�7���}VhKz����P�֮]��@��t��%���'�����5��o
=�5���i	�_u���PaS)��c�����;;;|a �;�&�@ ��O}�S����|w���b�V%�BT�P�0єp��PBVB+�'II���Ɛ��p*�P���'@�;�/Ĵ�H���Q��9�Je�����@,����yVE^�&y6Y~Ҋc�E`]�I4W��8=UW�x����@�gx뾚�v�'ZNjY�. �!�MTǒ3��;�·R�>����{��)Q]�J�:���	?D{��V,���yq�c˹����c�'�k^=�GN=h�K�^��z>�jmE��AQ!/��$�9�Ƹ؆�@�?p{�.\��B����?]S���>�>t�,��9ȗJ�t*�<hK��o����cB1�f�~�kV,g-�MIF/�a����;�vXDT�r�Lf���|:�쳝n�)�8	�j����P)8Y耇��:�
�m�}�}+���%s�<� R�x%�(>����Gs]=�"������tc���6lp��:{�E+��*���=���q'�^�0)p�gfM���;�Qk�[`C�a�H���`1T��o�����$��������;�$K
��X��O�AEO|K��z�~����y�B�}	ʕ�=���x��9a�u��N���s����~��۶�p��k���7
=�l��Z�ڏ9�h���WY��édS�`۶l�%K���֯[W�+���	�og�=Ϟs�qf�഑FF	g&P ?^��� ��b�U&??L_��|��\�S%P��]W��fϱ*���<�Ѱ1���}wa�h��� پ8���Kt�������AQ�SY2�c-V���~��� �.�v7cރ�NxQ]{��㋢Ě�'A���)�/F��ͧ?��\P��}R�.�)'i;�G�]T�:��3�K�����T�Q�W��(�/�fmA�~������;v�w�̛7�#���k/��^z���O^lV�X&]�'�\b�V���Զwo��`����{��v�igء�fCŲA��w�u���e���.���Pxw3�VC�c�:ʮ|߻�R�l�҂%[�~����{<�'�	�#^,��P���*6�������rV�~�eJ��� Ŏ?�|(�a���.�Q���h�8�����Ƅ;��,�����Ak��׿�NQ�nc��o��h�_c�@��;�ck�x�V�_�-�-V������>h�$�)}op�Ҁ�����:'%p@\8��'�Ē��西�ۿUVk���4x9dꣵ�e��4*ψ����x�b����ݲ�#��+�^�w�(B����A䟀�j��Wi s��W;ː��l������ۭT���N�J�N����vX��������3gz�2�/}�Z�0��8�7�\�](�yS�'ڬ�=�������:�+���G�\�f[6��m۶��Ѐ���&��d�;z�ڂd    IDAT��3`���]����ɇ�����!M�@&��w��Zil���\��_���9�D�Q�5
�=tl� #4�$q���}Ќ�Iʂ�F�_ ���}����[�h7���z?�񖦪��
9m�c�pH8�.ມ}�M�7�_�'
��E�ٗ���z�s;p��g��1s�L����.�3}b_M;k�s��wQ/�۟�2�4j|"������]���wgw�}�7jU*�? �/�B(�.������3U+�6ԷնlXc+V.��[^�D��l6o����y�����\iO��x?�������:���]��bw���f�_K��G�9�>�����@�M����n��.��� ֮Ya۷o�\��:�]�u�[�n�Y���o��N8Ů��
7�]�Z _� my�ƍ��H�yի^� �{*zB��g����*}��z�ȗ�ǚd��T_ ��
�����w6 �Ɔ��;���X�o��}H����w�+�BY�� T�h��rG]+����D�z�Nq��G?�dAU�P�E��u��FT�	�ڇ��Z��������o�AH�r=�&��g��%�g̘�5���|ͺ#T�dAA��X8c)��	��ՙ�O-�AC#�3FPP#3���07�&NX4&�q����d"b"Q.	J�F�^�`��@7�s1�xM��#q�Q�iA��޻����WOq(��k�jY���t�W_���<��>�rP�x�Y��M�Jc�����׭5~�ayy�ik��wW�o�˫͇��7�1�w�W�A���u�Ŏ-M(�i��H���<d��u�d���_�5eʯb��݂?�燆�������M7�p�|���<������Gc�MC�G��9f7L4Ti6|LPg�Ix�f����QGO�- ?�E����8Ё�<�P54 {��G��ի�Xx��J��^fF
�;�?��?}�o���Z~����[���Y�%��:�d�fu䘳>p���� T�8w�~0J.@�9h"�S���"X�6�M�EO�%
ȋ�"@1q���yꩧl �@u��$��3 ��/�Iu<=�("��RC����0�a'ث.��0����7W��>5f}çf�A�������~����ֽo�����bQ[�ߚ:��-��K��<�Lq���/2ш1�]e�������cL<�l>��cӴe�Ow�+LӖ6��ǟ����yo�f3��/��.���0l*�@J����ۇKI:"`y��[-=|�p3c������8���,m�S���R�A�C�台�.����JM7�dG���k]�G����g&���M�TI!�"�'��-�.�5� _un��<
q�|�X�d���Y� �|����_wQ>�f+�y�ր{��,��^ u��M56����9r�5 �V���QG�6���}�|P�.�$a�zM�ii��-M���%n~>w����kk���^�j���g[�IS&��m�$�����u�Af楗������d=�����<�$����47��`h(j�������ΐ���Ō8� ��N��\s�]t4�ܹs-/�;L�>�Eê��&��c�)�:@P����\௳ v�
�l�����MK��ϢH*��1��m%�FA�����V����hH��	2�~�Q�Z]Z��a�����~��t���C�˳᧒8�X��2y�9�G���;{Z�s4�C��|��]��3G�=���>f�wM{'����6�xȼ������N�HF̜��7Ѳ*Ӵ��zZ�Ye�?��UԖ��)S��/��P���G�0�~t�ikm6}*#�ŏ��i���f��LssS�(��ټ��ԯ�Ĵ�yf]}�w�?��*�}p�(��h��1cl��,����F�0dlD5�Rj�
Tz�i�/ �2�0Ȳ
��eec�0d|�,l
�y���}7�ߵ����Oh��;��Ϻ�R1�}�]̅hy�<X�Z��]@6S�Em�C`��N��@_���&�y�1��c�W��۾� ����Ƽ��-�67��_z�x�P3`@�z�*�mNUl�������۫L$��l�3�c�8�_L�>5�ݕ������?>h��/Z�����s�zZΟl�2���!f�W�f�;oϴ����+�j'�j~Sf������6��Έ9���e��T�e~'�kN�'5��xW�/]��*e(��\bU"��r��)p.���
��B�jN=�T�{饗� ����L�w�cU�?�%��^��N�F���_)��.\h���gk���m�R5�Kɳu��s���=7���+��Wz-s��o��k;v��������%ւR�<���iv��u��0��m:y[{��:&u6���'����]mZ[�滧�iFr����k���^��C�t�a�Ǉ|Amm�}E���LY�5����������ϛ��C�d�;[�����7�3ﾻ�������ܞ����io��ƦN3쀃�q�Oܦ/��Y��<��ݨT2rF���*
c��	E--�=��rnfDO�?�������W���(��{l�Z��(�02
�10 #
��5R�]�$'I����V ��G�=���v?`��;Nl���nO�
	��||,g/�g���b��b?ślX��Gٲ�Q�jAk
2���V�����u+͇~`�;�MUE�54�imQ��xɈY���f���jL��l�����y����r����Wjݱ�/Z�h�=���'?�;3�Ӷ��:�/�O7t�����g>��`ֽ�����?���z��N�
E��Qc̸/kF|�M�b��T����c�*Iכ�'k%�e �/!S��Z�͛2�}��kv����g`������m����ݢ�l��a�_Q�����R��B�?�F~?Z.�>���2(���X��(Y�
����qXQo��,�G��œ��>���Q����I��)�FԨj3x�D���7&�n�Z���_�����^5��wXs��:ZU��|��c��8ҔU��:���j���{MWW�Z���2h�E���w#�?�;=��O"x�3<�\p�~��6SQI5/�.v���&[�a��>��4π�M(L�0����8}6���S�G)�Hq#�p�|�@_���������y���!�s��P�}uV��J�T���ϗk����@���J�
HRTUc^�o	��S��8ܞ��M��U6�/�`S�|jW@}��/��v����Z,0�o2�ԟ����~ �?cٝW�-�L�K��U� P*R�M`�ޢ�T$�B55�S���Y�<� ˥I�$ݓ�l�w�3��N22��0~"}er��*󅹄��ء�m�Y�V�N���$9=�Z!�x��}��+�@�t��d��P晲s�ռ��u��4�4���I���|����oжй7�p�Ut�r�<yW�T�Ϝ��Czx�J:��x|���wW���B!�|�!>������U���o[ϊq�zy��4x��ŋ�Ut�����EA�Sy����T��iXm~��L�l(����k�͙��A8�� nZҲxO?���JQlmb��ֳ��ci۾(�d� o] +��o�l�w�y�n82����¸d�Ӧ�	 �߷��4�8Nm>�	��N�� �%����Lj��	��1Gw��{��ލ��� ��\�YʖM+�W��������)���.��gP(l�p�m�ؼiQ��ś3^��s�̖R��e� �|�?���i�(i�.G
�"< [�3�Ea�1�ָ [���@V�1'F�t�_����A��}��-��J�=�5/R��Q�F�8cE��9��T�=k��>�2{Q���x����I��}��r�`/
��!7_2�Z�Ƚ�KH'�I	�=��y�P��u��9)e>�{)л��@3n�eW���d{y^29dА鵵�w�O�2��Xl�iYi���^r�%i�P���2�u��p�b&GY�dA�B#+��E>���m M�g!N���D�p_���{�9��]ֆ�g����V��:�'VY���o��;����,O&���%o�k��l[��WXA����[o5����=�@�a	o��
�@���)�٤,X'Z:c�1mf��OA-Oϥ6���U�/`�����R����n�=2!0���f������<�J����?� �?�ܒ��u?���+��s<2���;��sm!# i��3�5���� BN~5�����IgO������H����)����d�k�0�k���y�f���4L�N�b-�Ħlz~�Y޶�8�:s�J�3g���@>���yF}�����K?��/�j`
Ɣ��xd���<�U��~;>�	�i��HnZ�<d����u�.>�8��b����2�m(ֵ�N�,~iu*��,"`ON?�}�m,hr�9T�ŕe�=%�,�[\"�c��h6n1�Bl*�q��������m2��ҳO�4�o斲�mO��
�;u
����S�>m��WUT����y��l&)-�k���x��h���r�=�	�]*�g����q����7�^��\��Qq��ѥ�v�`�x��z�H�\����SbN @��w_R�Re�} 2d�,�=�.�(�~���chqrޙg��>7Z�>K\�b�-�1�Ϥ�d���[6����c2��s�O��g��{}{�F)ɪ�QCCq*#@ԩ�J~b����w�� pƃGKJ7��Fź�]�}������C�e
Ƙ3)>�xP d��ٯ(�[/Y���d�Ew�O��(��N6�P��&�_ZWՋ�����4��>�$��92a ���
S�xJ���j�An�� (
E�k�IG�*j�T	cM ���u���J�rS0ڂN"nA�GQ����d|x"<'9�|�R۸�@UHV��R�6������*�Y��&��
�G�bL��8����]�Ck!��뤸v%��'�LjL�����di�&s�����҆��|����7�W<+� ���E7OR}�1�wJpd� �6m���3-��d	���'�p���/Y�ʣWF�֒�g�jf(�M��?8��,���3�z�V�T�2�}O��`��KT{�q�x�������^a_��`�^c�6U��Ŀ�E�fƈh_�oK��simm����)S�b��og�d�Xx-� �u�]Nյ�e�sf�YH�G��ʱT����D\�xg�ϱ�\���?��u��a{k��`|?���|��M���?�����pc��bG/rL���	@]�������������B���y�~ �>�:[�L���}{��~}}�H
R���񂠜Di���������"�2t�;�ȋ���Yw����nv����3�N��q���F@F�*��z(}_YW�||�Z��|?^�&t�,X))�����:�w��7X�^s�g��W�j�	䛗xz�${�1��Dɸq %> ��)) "�^Jo������/E��3�%Ydb�0�k֬�^s X�c.�,���7M5)�[ލp@^�"�H{^�\�EJ�>��-�������ű��)��_���@�)��N.g,�ׂi)3A��I�
�[�wJ�k�
tt��o}%ҁ%��r�c9� �Ud,���J�g��R XԎ��x|��tM�����/ZŢ͐���O���>���
��e�5�@���f���l�o���<3|�a�2���gPX��Z�?�Q��8k���ڂ�9����z�QGٸ��5�*��}tϋ҆:ԚBy�(AY��R�2p�K � |�M��K<��ISK����r�
�?�D�7�H�~�<���=��+�����9k��e}\�'��ε��KE�6��c��갺y�|])��xc�l<�ﴷ��(�[�F:��N����b���g~?����Am?s���a�R4�.nHaK!
oDm2���d e�=�Sy�:s�E�*>�2��X�qj6�( ��L����ܝ8�dIZ,�A��U�h)��7�{��J��od�5�CX ���{ �@��թB.m�*�Y?�ļ���nu8d�w6��!!�6c�!��象� �x"����������,}ι��=����$_���e+�U��`3纲A�lN?�ck�[��c���UJ������������V��D� J�C �~D��PV�A�+D`��3Go�����!N|S�f��D��p�}Cn>�$0��(*�/Y�X��/Xʌ᪟α�*'����d��k��"� ���������s.M+c�k�RgϞ�ND`O�	�-ݚ��d^dy���Y9��h<cP���衇ڸ�G���R%�̢.?�Y���\cEϡl#)���Z���amm�m%�O�����d�?�kd �X��d[ @���� ��ȹ��z:��H�:�`�m(��Q�6֩
L ��+Ț�Z6�F��~b���2b�� d_�m�@�����o�_)����Y	xc��I ������Y�� .:��� i��Rb�����X۠5b�?�я�gB�(
O)�xU�.2$\�����s�A@A2_o��Ft\����͂s<����{sv4��1��O ���� ��/À7��IW՜s��f���|�i^ޡ�͟k�H�C�"�,zf�����]��+Gm�0�JBI
�ˀ�U2��}��naݭ%����_�?V,��SD����
�m�`
�@�2��7����s�)w�7%%e��r�-�2"�!P�����L�����Oa�����?c����k���8�kg���O�1,�Q�F���41"����ǈ@�g��W2�I���\?�D�Ld��Vy�J]���|3>y��_��k�I]�O�N�VLbW���<��kkko):�<e�c�����h�]�0;���Y�JU�u8F\m7G�;�*�{e)�9e��9l�N2��;�;,�s@�Ԁ:Ԅ�����[+?�����9Wm���l��--�������Y��?��mV�G����W�})�".!�������H$}�D�'N�'�W���qO�X�7_�����}�`�h���В{����ߕG)�P�W4����7{��1�}�����̪[�h^с����o�&���O6�w�'PKJ��q�A����L�/ik��A�?�?����4���	 �^�������F��ˣ�>�\q���anPrk 7���	����s 	����K\5��B�?�r.�$�W@� .� �,(�ݦ8�b>�d�'{�TfёPrx-J��	�fƸ�3;�������\�����(�Cr,��Y`C�� ��|Emm��%���h,#,������
*+�$|�ff�*���m"~�}6ΟTO����(`� �7�'=��C���( ���PN��p}��e��{���x��,��Iٜ�����?�NcA2�|i��Q`�!��CB�3$艵��@�9c ނ|)��A�}��'�M�m(EdIVv�\��v�.���)��w.�_��x�����(h+�'S��d���Ʒ�ͮ[TwS�P��g��ם���5bQ��[���& ˆ<���m��
oد���dc 초����-��!(�!Ç��j��T;2������g�W|�8X�>A�6�_�	�����	Z�fX��z
w&�KcA�'���R�$�
���^
��"�f��W�&�C��^�_5��,�w7#&׶앩���Q�x��񳁿��w����*~W��(�ނ����S&�6�b�?�>�( ��<k,,�P�Kr	�6�r�*/I%�|h@��*<�N�Y4�8)u�M��1��M)\+�%��_�J������@�o	�}P͕��Z��1!�MX���?��r}֚���Ɂ�'�/y�Q�ɋ葇ӅK�c�C�4oi��#d�'�T�jŐK��ݲ�1n�I�t-�\��˂��*�E��mo�zO�[��?)��CO'qw��;�_�� �y��6���m�6�v���KdEʢ=��al����w��%ݓ� R���,.�
K���'e����w�%�{˟N<�B�?�?���rD$�Z6`���`i�    IDAT\j�'���@J������@ܢC��1��P.j{�ߩ ���s�1��d\1 ��y�.��<���������ɤx��D9�j�He��.R�ʣ���Ӥ��Naw��z"�-j���w�9��������:X�8�^X�p��9V/	�@��ķ�M��|�K/1���;����{��M/��\�2>�_U��L����](	��9�\h���� ���-rÒ�(K=d ���v��W^wwy�=ɔ���{s����3�.�e���R��t% ����yE:F$��y���/���x��������Yg���/�˳�7z�@^:�2���q�SEn�<�WM�,�'�|�ƕtɹ
����E�6��M�8hGɂ����ރ�Ҹ�]�]�y:�2��E�a���)Si�5��
�_@Z՗�'mjDux�(�Bȱ�iŠ�Mq��բ@-�y^ �9�?�n @W]lF5�S/��x�0��òǺc,�r+���/@�kh� �����k��w�A�(z������]EQ��/pI�d�駯yU]�LGb.s�*	? �,B㩫+S��52R
�x�z�W��ǖ&t[0p=�} i��B�P(�G� �T�r����}������9�w�F��Y�ъ�zRT�5j�o�(V�+<���0��������ŗ�?iꔇb����S�?̓��`�=A���b8u�+��T� -B(���-��O��=��-<?����<��s����K��d�;�?@��/}Ɏ�!��q�3�=\P��ML�7���;�$�K��d{�m�l3CRV?���~�^
@�� ��?�{���ώ�K�S�bs.P�okB�/T~r�F��5u���]d/�~��;�3�?��24ħ�� �mj��R.R&:�:�X{C�=�<��C:]L��n :��>�߿�GO=�D�w�<e��i�5�!��)��V:�
P#����\RH���XHV���Xx+V�H��U.����	����`s2ר���sp�ƹV�I�5���a�A?���h�"[�K��P��#&o;�KV��)���y��S#�<��؊����c�  (�����l�[)��v�gw����u+b}�I����#�ܐMƩy��� pU��|'ʜ@$4�:X� ��c� �(2��3BYI�!P=('��w����'�H�v,͚�{f���O8�������ŏ_?��S���5�Â��v-��@3�� K)�XH_��K��B��*vt�M��f`#�7���j�q�]�p �i)�����e~^�� Y]�8��a�Gi�P3:>�s��w[AwG��T�BQ���Z���P�� �m%�_�M���m1^x�U��T��ۄK�/V�w���a�J�����j�u��\�C����:~�Oz����O�|�^ �뮻μ����j��?��F���;ڲ��i�9�5�a�o�
���{�N�U����S���"�V9D�v���1"`|]��;����g^�0����|�]����O�')�vO��Y���*�d#�	A�{6  Ϧ@�-�ʝW{�̞��VIc.h"��s�Il:�uF0o���ҍ�Ld|6^p�9���`vu���#��5bx'��k�eA��I!�݄�/��T��\p�����r� P���S
�>�\|�V�*O9h� ����i���h g.�I�k�	�gm����?�Mx�4�|��Nu�d�-|��U�(/Q�Ɍb���.����j�����l=����x�s��a>�У�)B�r[cc�=�~XX�x(����mm����aWf�,���7��T<�VV�{������8�b���ӛU�� ���X��lB62uӗꇱ1F�1��6�!���(*p��#�1�?���R��ݼ��<��)N�˟��g�.���,D�e<sQ�r��$)�C�s���{�N�H .OS�G� �oϝG�U���2��N[)-Q4���߅|�{d\j�#ߜ ����I���]9�U.�x�u���u���o\��-���L�n��ƫ�T�OgJD�v#!�X�X�:��M�S>����tK7��0!��'���@�?�B}�y��C۸��5�Rg�jL��;����+} �j����Ac�Z�j�Z�|k8���-�K��6P1�?����0?�?��%�-M����8�Y2&o��e��d��1l|��	��t�WkKO(*�m�>�g�)��ؖ�Ke~rO�_^��+Y��TRyԒa�0�H���>���[����4�/N�k��������oO���'�3m~��!�m����K��4�":(�'V��$]�]s�VѲ�]�K�#��Apw�M��`���i� ��z��d��]#���Wq�֦n��.�W'11�dz�y��f,�yF2MHC$3��J|�Q�TO8��LJ�J�eZ�C�馛�x�����9Y��b1�7�с�2����x~h}WZv�er�g�X�(`e6�5�<gbܬ��;���^����w���a��3>,h�V�#{���O�~���z477x�7�y�O��7��Ͽ���^_������W���Now�Vs���Pv9V�<��5�  ��'A`0��O�P��݁��YY��=�!��( �� :�Qx(�8������K'�i��o(�e��pjn~
��W�=�%����g��y���`���yꮲ�>��������ᕒ�C\�s�Y���1�8Lf�ܹ�������J����&g��w�1�ͳ�<�[�w�ڢ��|�G|������l����=��]s�����ٰ�e���8d�����)k$},A>� �H��f\46Sa�t��`�ɂE�͘1���~hSr�� ]�E�qh�[Z2�0�^,h�rt=�B �����O�Q����k��?���y�I�ĲG��ƿ�� �W���Jnh��}d��k�i�X�6��mW�|D%�g�d˟uW�+��θ
����e7Ͻi�	�����9��˗G������۾� ��"���D覻;�+�(>�wQ�*+Y@'�7����lyv���H�� �A"*�`����)� ���;��������aEqo
��P��>H�$�"CF']1&�
�����߰�I���u�.�ÒgO�g.)�c�PH�A� J���w������$���o[o�އ�=�3c`Ȏ��x����.Yzaw���3��(��O�x����Y��P�]*�W��-vw�����С�d`(8���Im(�_�)$��͟6	��un��RN����c����= +�-���q= �L��Y�����KA�����Һ@ֿ{���f���8ԅ�o>�Y�FoZy�V�?��5'�S�H����'D�
�WZ�^$��?xg0g�l��T�2��ֶ�	��y��=[���5׌[��s�Ps�ҽ2b�Ӽk����_i�n_ײW���b�\|�S�gf]�gm<�,�Ϳ��J������a�Pm�p�B[��D�?ܿ2F\�E�|ƯϺq(� �5k�=xE�\�	TP,��]/��C� ߮'�{*� F��d�`TA��8���6̤%sp
��<M� 
��ۓ�}���7��Omʭd��.���rS�Y����7/�q�)�?㌕E�<��c�}��~S�J@���}������XG��4Qt�jS��|�3��<7cb������%�����8M�Hl,��*�����Z��w?�Z�����d4�����¤/�I��yEQ��"Њ�̳g�>n�:�Qv��?�?@��!������Vz+nB�k����ϧ� 뎼�P9���s�I���7��������@��ͦ�~e2�s��o�{�-�A�����ڴ����sX��R?p�z0ϻ����`��"q`!���Q
�R�5�LlO���SdD�/Y�
�a	`j��P�?�x�Ny������#e��w�ːB�'=� N]�tU~RYK���eZ�x����?�wPH�h���T�>�ޟ������/c�R�������<��axfd<�_�}��˵����q��յ�k��o�qyу]]ݨy��-����6 �pQa��%`^�޽�孱���&��f���t?F!�k�Me͕5!J�9���LOr������ٹs*��wS%L(�2Zb�����9p�pǀ����Q$V>Y.��
��J �'#��cUc�B��=�>3�a�ųJy���ݺ㡭6�N��3�����g�bW�G0n(�y�7Y���(�"�L�//]�9�O������~H��+
�2x�Iz~�p(l�xZV����]�.�P�����z����s���:l��t��m�1�c}Y+�*�tXŠhT�{dUQ�-���lsR����~�UH�b�T�j�\�ϧ�rʧE�L��i��[�z���x|�N��F�
���%m.ޚ�G>7�c[��[����'�! �r����>N�K�\��75nN��"�)�&�w7�����E_��<U�r����`�*A�� ����'U�X�|�@������J�T1���Bʏ;ܟ�S��HhO���<�h�J_Ei��g�� �')�/���y�駶i얹�p�s�J����!�#wj�)t7��w����m�������-P�ޙ����
��a_�l��+��<3
�y�M���O���ȅ��HH(�\tw/��XEvvvn3f��{��/Z��*ڇ�_�`�~,�;O?Myy�; ��E�v �F�:�r�7�Y��>xܸq铓�LP�tEU��˃E(�Q��m�UQ����L�|��L�cu,_�Zuڤrְq�f���yq���.��Kyq/�	J�MN����g�B�j�\/���t��m�V�*\h�p-v<z�C��l�%p銟0^�}��Ȋ<��s��3�ِE��SOn���sJ�?��/�0�̧*�W�[�gf�Y�&��-CF5̽���ho�b�ʬ� ����q �]�_�N�S+y��DQzmy?��dXN���k�O���O<����\~��ǿ��˿�ӧ�H{�meEZ�܉��s7C!�����r]^�,0�!��e�a�;6����Ea��Wm~��_Z^V�"�Ue~[]������TAO�M�>��yYm���㓲�d]���D҂?�̼(��!&`ѽ�,�^�	�wQI���O��z�(p͸�QQ�'��L)@�O�QAA�>���m�E�06�g���4ߋB�Y�lN�G�b�#c(��z����`�R�G"w�� \zO�\4�s_��%���}�q M���p����_��| �����U�<���^ߵG��Rm���rV�?��y���)h�����'�|mCC�%����9�J�]��K�4��D�ȍg��:�hk7��~�3fL�e�F�eVL������}��g-��� ��<w�)�9(gS��~7��sdZ��m9� ~�6(�Ϻs$��C�v@�����/����(%'�r�H
Yi�Fۙ�5'|ʊ�'2�zi���~P|tO�z�q+;H�,E!X�����/�} 8r�a3�%�Sͭ�S���_~W�T��p�G4��h+���kC���[�-m��ȋ�^d8�.�K+|ݏ�j��.�3k�Y}�n�<�ӯ_����_��#��ܓ�/:�gRx��!,��L&OE�宥�����=Y�\׈��e��a�6iA;��@����<����"j�,�_֢��I�ϊ?tw��y^�Τ�D{$y��M��pĔWT��]��d�+����w�G���a�1?�ݑ�v�$4�X�:V��x�_P�T�P��QO(��K�R>��9�oX�dĐ+O!�㓬��c�+ݏϋ�p��֓�c�/Y�����z��B!�G&�%=�C�א	��UUU՞�<���:
U$*�=�]�s!kY�e\娹Ҙdd�������s�(�C{j,'�A���sT4/��Mw�W �L�%��m�ng�J�gȶB����%���W]u�'N���^E	�����_?lٲe�&���P(�E�Z(�mƠ	-��|�����
�d��
���cҜp�rQv|7����wb���-mQ%����/@K��*+��s�Y�9bd,�G:;;�^�y�U�!Qc�6lذ���/ZB����,:ml�'�S�G@�^�������ŊP��6Q^����B���M�Pn4�#�5BqṸ���nZ�ƪ{�l+V�X���}�z��6TVVvvvv&����x�kkk�.qsss��7�<�����D"1�ϩ�R%N6�;ǢQXGY����E\/%�idz�?��}�dp���ʢ��mŕ	'�Tb���;]z����P�+���TC�ВiӦM?������E�L��W_}����vk8��#�b�Kg�t�����u��7+@R���h�vԑ㶩���=l e�P����Ӡi���.g�qh=C�����)P�(-��O���֯|�+����y���jmm}���	�*|r=9�f\�R:.5���)��,���<{�g]�s)և�9����Ҧ1�J�m��u��ׯ���c��3��,Y����n�<�L^TQQ1P��F@�m�P�R)))�LP����nR>�����^����I��C�6�#�S��{K���!X��V����>�Ogg��&M�����/;r��&j�̙_x��7~���|Ruuu9�� �+���L�uG&�7�u9J崓�uhS#c�y�\�6 ƺéM���V�����ZX�x�O��o��/�~�ĉ�͛�yPvwwvv� q�xpV�y�mv�����92
`� `}}��	&��\���5���/f���\�D�)���K�i��5k����WJ�QG�{b�����I�V�y���	<>eE�{��vw�()Ŷx^e7��ʮ�3%N#E�꥕����&L��ùs�Ο��H����Y�f�O�YUU%��!(�rPQ��Ke��=hs�|)v�J��pD'%���~6S���
���s�euf~�P��VvGJ�mPS�ȕ����1��a��{�wP"�x���k��/�uQ@o�fv����R�t�u�]���N8aNO���g���[n���h����d�E��Efܽ o*����\��mI5ֳ�AEe��� �:�*���������'��(9A�O*J՛H$:��˞�������:�����&��;o��§gE�E�0�:g��M 4�S���{�.gs(Sg�j�i�e���E�p�����M����8_�?���W�"�HcMM��ٳg_s��Gg��S���1���NS%(��L��<=N8�閿K��A�,׭[��c�=����|�w�q��yvuuUD��#cU��������i�lRY�/���˭�p���|�S�Ac���x�{|�ғrPFolll8p�G'k�܋/�8�>�5��;����O��������G�WS3`BWWW�F\�@�|a�I�m�P�����o.�W.�v  �O�}D�d)��H��~��UJ��Xuu����}͸q��s	��yh�%�+�1�(h+�_ ��"sn ���[���	A�$_��*풿�8��L�0�P(�p�'|����Λ7�Ɩ���*��?Q�W+N�o\HAle�Q���ԙk �2ʌ�� �έ�����O���gd�RJ!������C�wڕ�>sҨ�:�z	����n��sK�~�g�S*+*noo��!J$H��6o>��g�N����~�K�2H[�X��&+����t_��� p"[���i�a��[��kN:餜TOj\�c�<�+̯,~Q?���xBA��~o�_���;>7�@����q��{�8��C�P���:��˗W�r�-��dӧ�VTT�+�\oS
 �s��Bge	+�!��������A�G�ic�{����lR�*ڔկ،�&����k��j���5gΜ���^k�&{�=.���#V�Z������-+UQQQ#�I�-�Lv���l�&�|7�M�e�g8Qy6B��>�΂�$�������o��7��>�z���d2�`8>��� �G֒� ˾'߷'_�&��A/)�mݸq��cǎ�rG-�ǲe����_ߵ���*p��.�+��̜�H  �IDATy�C�T���>��/�V�	$v��Lr��^A�A�	��h9� ��ۦ��������:�����g!���=�͟��g���u���S�x_����D�	�BeA�Y��=����$�t56�/碌��L�l�dM�B����S>�+�r
��M&�=u�W���O��ӹظq�QMMM����k����,)
�h��+(�#�z{���9��3f�V9�1�S�zÆ�ǎ{��X�����ȧ�x<>����wSi��1�}�qf� �A�c.�WO&{-�4�S�D�o���}_�-?m�p�)2%����Æ/=dԨe�_}������%�߁�������y�o�f�ڣ=/1���r0��1������G[_���m�c������X��l-�d�+�F)���(�!zuvt�C�Y��b�!���dk�,GnL(�[�!i4e���I�?o���ow��ߞ����[��0&��x޿W��{�ҥKw(?��������YC��h�H��СC����&�Tjoo�ڰaC���2���E��]�,K�·��gw�}���9C�2g��i�������p+	�{�����[B��F��^nhhxvܸq�������˗W�����4}��}C�P�"��}�z���^YY�d!C���}��uo���߳�dS"��������(e���3{^��8����Ic�e��m7���D"������5;�Õ�}]���m��n���Vw�X���i�<�-�յ%�%�G��F�<��G���СC?�6mZS>k���R��Ʋǽ�dɒ����������6m����N$�
��D8��ɤ�,�3&	A�d�/[�掻�q�{���F��x���a��q@�1i<�Θ4.~2N���O~�߾��"a�ya/�¡d(i��ԘӲ��1&�������pg(jO$M�H���΍w�}�_�������w�jjjD�����Ӳ��pWWW����-�d�-5���ye�%�ɴ��L/0�LF��p��<����T�B!�3�L�<��o��S���z�k����9��K`�����RH3�]��u���d2�Qc�t��y�
��P�q'��L&�{�GH�1���J$�Ϝ�e4jMd��:��h[(�t����9s����px�>}jR�r�|��i��~�`���/o�{����>ӽ_����R�;]�lV�<�8�dKE}��P�}:��%�:]��ʪ_���TD������ͻ��]�0s�ѿ'.�{��k����m�lI�w��Qm���*/-��'X<��j��/�Lߗ�~N�Iw��~u����Q�G֩.�~NU�6t��Fc����q���K<"y���!��ˉ��g2ټ�OJLI[`��j���A����mP�C����X��9�?���cfAt��S�b�b��_)��%��i@k���1O=$���&,� ��~.�� PK   DU�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   DU�X(	��I�  &�  /   images/b4edf89d-5842-4488-bd77-04cd2da60bcf.png|�uP[�6�'8Žhq'8�R�����=@��ŋS�xq��bŝ ���M���~�����̙̜9g/����<k���"��M�  p�߼�  �P䵂���#����Â��w �^���Oe^ � �W/�<3�31Ԟ�]ݷ�=8��36�X�g���r6��de��O�ɡ'z�����ל���f1�.��
���E��q�\�ѡV����?�m�_���\��g6J"J �o��x�z(��+��	�p�����������訯at��:�����<3*�����0���B��U>~?9�%�# ]["2�c;�^���5��6��n�Ba�|��A���1(h�]�I����qaAbO4����^��7=Bcuv�&ۑY(�zL�$���\úҋފ����2/i�K,�>�����-���р;�����(m^�@@ c�?������8����`9F/W� g�~��se0���A�
���m��� (m�8)���||�o0]M1�_UZ�{dD�����p�;��cy�O��&2Ouc�k}�r��A�F~�s-p
B�� �oO���j߈F2�1�b���>q�i<A��N��ZC��7;�FE��⇕h����š�#� .�6����s���x=(�r{ǽ�-�P��
k��������>��k��e�ܔR�%F����+*
��0�Ȟ<W�琍��E,nsc�r'0]���^p��d��mvL-W��+'D5�W����3�"�H����O9�H�$:�qw2�-Sl��b�B[����E�LNO�����h�WÅ}Ӟ�vL��=:v|�k��������II$����_Hk�O�+�Gh{�_e�������i:>e��\�+4J��+��,�f�Gr,Xa�.���z;;u�/��4<:t�[���T�����n#5�aUN�ι0����B� WW��qqq�l��
T�󘬆�&:��X�꼁���9b���T6�Wts8}F�/v�A��X��У˃7�s��87w�.��L��Y! �`��f�PO,�/����L	�s�˦�Z3ӌ�w�=�F^�Z�yX�g<��ɱ���!�+9F1z�"�I�8���M�� \���
5��C��,��ÆÓ��w���<�_?����S���~S1
-�ΈH�Bw��R������7��,�s[Z��:�0K@i�bb��u�CG�1���(B8C�#���|��BE���:��X���ڔF����r��� ���'	�"���.W݋	գ����g�����$�'qs-��#%�p��^��h��C,��(���!�][�z���J�[3	��6���vʑ�\�)��=����w����8���'��m�C������B������D�8L�@B����!o�n��!E� �nq���4���7lzzz����%�����o�����Q�e.|5݃$�}�r;� j�&[k�}���Z�Lw|:��iV�����;��������+23A\Ibc���~�9����~��40�l~5K|/y��e��X�K5}}���ɤ���{���b�45���|)���+�T�N*�JTO��R`L�������o}0NC�:-"5��n�rDd�|O7�s��أW�����u��z����u?�Ʉ�׃�C�Fv��&	��|���{:q/tS�����]�E-�j_hA�[#�G����Z��T�}.9Ͻ]\�Z<=�H�W��K�aE}��W`�-g�Ӌ7�P��`�P��fI��?�6Wkf6�e~7�
�/s��LW�{��J��kX�)����K�x�ֲ��$W&99yr/�&(��lhh�9������&g�c�+5�_SQ�@�Ҏ�u�NVu���-oPEj]�tL�=]^�T�Qu:lg�/�`~{շq Q1�B+��@�,�GFb.n
�Ӌg�JI��CW�AP���
T�ꥊ lI%�"��9���q���2Md�Q9�Ln��h�N��)_M s�U�q��z�z��җ�f;	)zU��I�<��>����ˮ�PPTH<�9�6�S�Q�a1٬R�����E�4
�1���y����~A����[� ��$b����|q�3QTBP�p-�g�	[�_ff�9:��^X���P�{c�`�$� S�˗��GA��=���&��y��csTc��2I��Vz��xUs�wg�(�h�ԗ�3r�K,�ON�o|���ߎyE�� �-�[��/�6qU���Ui���zag�/��x�u��:�)���7���O�4��H�� ��_o���*�f�gJ�	��'�v��ZOd�_pPP���З<!�����)���RŢ�bΘ�~��L��J�7������~�����9`�~�4�c��sx;��eǘ!��d	t�xC(v}����e7���7&$O�����{����H,���BA@E�\�e_LA�����m����P�'�v��Q����w��VL�`�A�U����=�t�H�Q��5t���MV�� h)�#��An�Q��h��YB��7kIh��V����[+��ދ�-���Je��~�T��TR5
��ձ�mYRb�����%?�y'����,LC%�(��F��ы!��m����C�+
�(<�w/�4^!���5�O�yI�����u.�v�yG�Ԣ�/K�]����/�4S��٨4���v�^��V�C�w��###���?��m�FJ��5��w�'f<j. Ӎw培��WU�*��8)h^]�L�StC d��7e���7%^�E^	�v[V�[x���;�+,�������l{å����s �%8:75=�͍���L�i�ozϏ~lbɯ�/� Dni��\��I�C�hġ4��L'�A�эZ��@�b�J%���/.�b콺}FJ�50H���5�1����-+�^oE�t	?��T��Ce@f��0��?M�֤z�,gGm�[�i��Z?w��4��B�d�Wj	[�v�u��y����@N���d���js���J�j���	�[����6�rc���T[����$ಓc1�w�h:b����*:�w�dg��0�ԏ]�<�^{�_|�3g6��#^6<J���b7(�F��Y��&6ev�-<����7
�Mו���)�[7ېa�Ҧ@��o�,��_F����ռcx^R�6u�'0M�%$�5�搕 0�Ć��Ļ.6��f��o�\RH�BZ|�����`���=&t�(}~���K��K6d�b!��8�<Rxf'XхJ�|��9��h�v��W���t5����T����}�����}	(��Ii��wR��(p�/�V����"{3���M��+;2D*p��TT;ו�M^ޠU�F�Cf�Zr3߈�Ӳ*&��}�_�+G(ۧ�0�߂�Hc\ r4(���uG㗝L(N�w>���F�D:��؋��ӛ�z�IN���̜�/]�W�&�'�!�~�� �W�o���c]�;8�Db	o?H�Tp}��'��8��{���"OI!4����_���'����Mg9��-�ѝ����Av�sxhwV�1�5'�5^���v�R�����\�ZW�J��_xdw���H������s.CaaT�C"�+��9H���p�����dT�p�J����q�X;��5��'��c�����mw�h�C�jKK��1�����ld���~��x~~��b��w;Tķ����V�Ë��[.�!%k�q�B��~�Qm�~�#gD��ѽ�`�`>,-�΢��r�@�6�����{�v����'��7��o)��GDt~�����ݬ/�&.!A&)ݸœ��|���g��W�w�)ł~g���P-�C"�h�_�P,��S`E)Ӕ������}L�����)z�ž�H��(����|*X�
��}О���N�w���FgҚq4����ɷ�P;Ko//uR�f�*A�P��W�5֣�J�J�3aϟH��t���,�c��b@'W�{�\��ٝ��IO���[�٪ђb:�����Z����A&���ք��N?�m��7y ��'=R�g|�*z:��e�d���B���Jt�\�5���|��V�$�^���p�n��p>[\;w���b�`�C�2&����s V�������!�%3okJ
�RF�M�����lU�~��. �Ϣq#u^��rONj��_�U?j\F�:9����+�6�.��Q�2�ѓU�����g�ѲZ�t,�|�{CfK(F�Q�Sе~�����,?�-�(�'|ΗT,`7;+m�̦��O����j��8)**�s�k�5C'��z���A�,�ZXZ6��
ܬ��9>�>ggϏ��z�@�0���1+�`�ZW|s���\���[5�8�XjqDhT�4� ϑ
b�W9��H�F�F���i�8
 ��VWӄ6tϛ�� e�b�� �-�T�ʦ��Ю��*T�pn�rqN��.R�)|O�B�0pg���CX`,}�m�������b���'�9�C�#��M z��_�N]��>�8���AK�b6o�	��KY4:,�\��҅����e7H�1h�xm�'��/�$�^ �ߜ^�w)۹��8`y�0��A�-g"\��7�P����r��OZ��b�P�b��̂
$�I���b
���9�d(y���QQ�������A��,��B"�C�q����fig�&�J�1b&bĻ�S���m.�{��Y�?�sZH+��}�����VPP@R�՗�(��	
 ��譴�{�]�o�Ч�(�W�;�cѯiO�j͂Q!�5���������;j&&�~�?U
KY}V$�����m��-�k<h�v�Y�5b��tP�����L\v�s�7� ����N���_�NNN�@O�1�T^s �	7h�뛫���/���뷰�]:ɔ �u�RK�'T@>=�S�6,R3�D��K+r��h9&5�1<���FFeB��[�1͝��-���g��i� ��f̡s&С�<��.�%K ����pm�#ݷ�7cYu�}�R��c;
���;��t|�~hw`��?	��LH��{#�S|#BpK+���䠟���}�Ԁ�G�&��<�ha��'1mz������c��PSa���=Ay�Q��=�<���N�R���i1�XR�شݠ��ӋTK�G�h�f��D'5�����vҏT���[I�\�gfcD\���e��*�8_�٬�G��ue�cr��:��C�t�*�Ă7��^��< �z��߿�UUU}=%��c��mk0b��vL��/��#�W[��S7��&�3/��T�&G�
�c��m��:R��Cb�M���2<_5��c mݹ��tQm4~|UP�̮�C1ք�lSh�6�Z�1�Z�6�瘻x0I��A�5��������s���T�m_D%�]z��?f��h�U#�꒒�����F�n�:)�i��� �Y�	�d��q��9-C�V�5Ԃ�����..tZ	4r�����c�#���'��!W�� �
C���2��2��<�50�"N�羹LUR�t��N1C�+Or��>��+��@�O�nF�/N9��ȩC�h`ˑ���ʎ��9��糎W��� !<X^[�6�С8��M�[�q.[j��	���7�!�
'�6��C�Ǳ�֩ۼh��q݊X����D���Dz�����#�(=�0*|�z�u|�VUj�о㥧u�%������SP`�{�D�B2��01qW3 ��5SV:Z��W��yы]��r���50[��A�A����ُFL�Iv��s���r���t$�A�2@���53C)A���lI
l<R�������ִ�;!J�ݲm�B��fe{�q'�`~���Y���︬����T���0�?!�o�8���������b�|�wq�Ɋ���~����c�;�'�o���dO�"(�pӎP�>�_���g�+�̈́���g��ZIm}?sDU�|�Hk5�brk���S/���<W��;������.%��ET1��l>E�I�v��DA��3���1y��x����T@��^�mt^z���0:�Vb��h��(�;P��]b��Vy��,�)伷�I�1�6y��IR�c�m`�� nSq��Ħ"ә�Z�;����"�&�9���7#X!�*�i���FOJ2(+�a��kp���Ȝl���)�H2d����$y3��xR���F�N��h�������k���p��̓�2?H�/�f��=�WS�̖A^�/~�6Z�6�Y�]W ��m��K��	F5�����Z��b�����X�Dm��'��Z=�;?>2Lp�ay͒Z �uɤ�m���f����i��Sȣ��Q� v��vf#�%{tI�����YQڰ���D(B��������o�^�Gw�Sh)���	��ި�O���Z�M����k�N�����@�`��;�cB05��SO�=�6��5�*5Y���(���8'ъ��@���l3����KL�E\��W��<�'Mdr��*x`d��@;b�NS||S~����U֦��x�m��u�%a������қC��R�-Q;�͡�pqJ2��L����Emj���sy���D���l�����zK�6�Z�]c�����Zy�ئv��i�,e��Q����ɠ�!�q�α_R:����^��v��{���W�ul���^~~I��&ϓ���>0\KAA2S� eu\{NIt����&L�����5,X�)_^N�����;�.����������5c�ލ]s�"��ȋ���-V꿚H�u?��j�?=p�����Ǝ�v�~���
ә�sdC �����w��\��=��`ѱ^��yG�]$MN ��7[P�v��_�n�NƂ.ā(S�<�Yn��@쉊v��MV��1>A�s
���8PvzY��W��b��t�^|2���|.�I�
e�]A�!�t��^�Q�N��]C���6�*h�6\k�z[;K��sPE��C������@1�?�ڨ��ī�x�.�HMl/k�����kQjĶ��H'e�I�@����q������]�;�X �ݒV��x��Oq?|�#��U��!�%�0�
i�����}�����Xx�����P��LX��S�\��cL�GEX#��w:��������t�_�������~���R��aZ�|�w RW��j�3�#��S�3zU�94_�k�ӛ�d����?⼢䑨�Ju��P��8O�l$�.G1�Ky=\R����t�
��dB�RA(���"4�Q�J��1�Kl]A������+��֯ʰۂ���y�Obb�9V8����K�V�_�S�.Z�r�w8�"
�VH���+r�n����9Qn/	sN�[�H�����Դ!-����5=���AL2!�� �t~J����ͨo��2n:���^lTd��9����j�N�Ę���.N��6ć�����x�Fl����H0}m�l)d˭B-2����j>i����八�0�{ukԾ 0�+���{����Ov��r2�.d��A}]�n�"s�n5%�l4�ǚV�+�6F@}�=�
Ȯ����=����R�g"b�5<2π�_����� ]5L�ژ�HȈ_�E|[˂	V#?� �]���|�f	m��Сu7�!���h�[)Z/OL�rn�� �4
�f�;���)���zg�C�ww� ���@P�<���t����,��eK�1���~)����5H��tMI��a������8g�=$ @&:o�o�6���1�/�`T�,�B��0�l��[x�
j�yz,���)2�5s߰����4g�:`#H�}7��Xf�?#��oRv���'�]���U`" ;�G�hic�O%�_�wq�M��]���T ��LI�,���c�%Z��jw�+�sDLU4������)���ɨ� g��s��[�*�s	�J��P�R3:�4��.n���fro�vB��~���w�����ov�6D�O�8ꀜ;��(���n����`�΀Uk#`��Ϝ��oAAA��>'k=�����F���+([+�s��lV�E֑�I9�#��]u��E	��z4^L��4
��xe�p�-��Ӓ�ɶq���}=��1�]��AO�^��ˤ��N�?��9��oqU���C��mGӳ��F�oҠ��~�v�m��~u0�"���6�e�kk��g��0���Y��������4��o�����W�3�����a:���c��+����"0�� �<���PGr-%	�b#!'�L ���jTf/�{+e\=�eM�xc� ��(DF7�8c����<���j���+T�F��T�H9��3"}���4����;�b�VZ��^bX��Ķ��e^��<������/	�Gt��w.�ܔ(p�=�b�Vo���uY##�;%�)0��7s��zH�{�e��G��o?8箭?5�(c@E��A��<a4�8K)�H��*8+��|�(6���A��O%�Tz���`��88J��� ���ٽ��f�;�aட��-f�W#��/K,���ۗ�Tн�Il4TUt�[�fA���������]k;�J.��|��҆�O:Wc��3�V<��YdG�P9c!��S��y��~)��_o�s��X"m��DX�����y?6�\a���9Xl����V����#�������/2����͖qt�D;�씶��Hwj��u,�wC.�5�a��)�#�G��Qz�G�kx^z��� �x�7�F�Vo��k�S���2D$�l&�)�|-,���<$O.VZS���[Ldd�E&�%z�yle��N�VY[pp����l�vn����'@���U �E+�g�g�	=����~�����2���uʜ�|�����p���[I�ӏ�P����Z��������������+���BB)XP���[�LӼ	bY����>AǠ�q���ٶ�tC���gtH;�4I�ם�
�x�$h)��ﾇu��bگv�v;|� -ظ|��.�h�@|.�Q10��bn�Z�Z��?�c)��������K�:&���|>�ʂ��Z��V	�Kȏp~�MD���8�`��4�ɰ�5�(��(�4J�����;Pm�`ab�8���� *ޔ?�b`S��_�2_�PC�Z�|d��L��\��n���1f67�D)�Z
�d��)�&���1,�j���~�{)��ݕ�n��m�69�I`JpʽF9ȷ��j2���]r���������~5�3�y��օ�w�C�T�������������߭�Z<O@�14���ŎK���G˭�� ӷª� 2v&��̽��\n	�����!��΂���F��ohWm���WDf2-�5���J9����,�U��z1�B�:����B�H����b���U�/�g�xq��S��-���9ү�,��_l��V�@�w�
����|�������ih��U���4T�ȁ��r�k�� j��!�G�R@6_]brbU3m�=`�&�i<>2����?��}%/<���zg0%]P�l~VC��W�ygT�iX�X���d4
�����w�)�����6%�����{ǯ�EEk�"�#�2%�� m<渥�����0�ס�7fv�d�#t/o٭di�@���j��x[BЛ�HX�>{���ܜ~\V�JB�O����4��cφ���;�o�@ϲ����q�d�'�];O�O�@��x�1.��I� ��˚O;���e'wW����%:xB��n���Zmoq��(zF��Y��S��1�݃h�Y���ۏv(-,�2���]�E�)�-�ٻ�������;n������K"����hv��2���O�xE�J_0�[�����R�� ��ҵD� jYJT��ZԨ;���=Ũr��J-���`Ѽ�.m�ω��F�jl^�k�߽ڻ�gA?a�o!�VB�ǌ��!�H��ĝ���RR�V���X�!�	>K�["�1ʋ�����Lʌ�)�v���c&PA�3�?m$8]��Ƌ��	�G����O���0���߼����T��~��P4�?����� L�����;?X��
\���,��1���2���r�l��_�,��2aFFγ���8�y#!1���R@��|��84�?�G1����2$O����1�oyW�c��Y*�q�����\ �Q�ְC��F���?#-����#.�ia�K�31VC�(MPi�
����d~�;��>�
j�f� ��VW�!�>����iVJ���EL����{� s�������ׄ����f]�tu�wɼ���2��C�L�%_��������{:���~X�l��

��8<#|#<�O`D�z����9n�� F��yN����`}������' B!�'�5�Z���x����-����+�𓮷YK߇��T��8\j�.�R�m�G���Q�fI�h��7�ڶָ�Ju�.��wr�q�E��>�f���P�;n�R'b�t��q�T1�n�M�S���D��x���W|s��(�ȅi���!�n�5쒨ק��T�XW!��٫�_Sb>��ד}6<�q��џc�ꃘ�t�y��
�,p�4�t�,{��X����A��-H�8e>X���?���%fߢ��F���3��y��7�WPFj���/��CR��� �����MF.۾�F�)��p����F����0��c^=K�����0��1�Y9��ǉ�sq�����]�׌�V(���|���?��cV�
]��}[�A��³�����5�9/}
+�O���J�0�
T�%��%����<΅��'�n�U��'��Y;Ѝi��vv	%���qZZ��*'��m6�6��»���&��&�^��OD=���^�=t�ѽ���ꋡ���.թn�:ϕ 8lG�׬/�C������N�liS�WM/��4�[-�ڲ2������=�$�'gozz'}��f����X���<w)/�$H�(�q1���맘)��X!�$�I����sh��g�b
'�*)��ɯ$b+nŎ�Do�z#]A�^Me,��Pf٩��sP����O�^�$�-P��,�b��p%EVZ�%3������%��]|�P��9�)\���"���g�sUz'��Ǜ�TD��#�X��,i�=����$' `��4��~_���;����'���o�)�p��=�Ju�Gכꦽ�L���QJ�t��Ϻ�W�T[$}�h��:\bG���fg�/Fy?��c�q��Լ"�bl�`���="�����ݟ/�E�Վ���>����=!��ާ8m�U��X��Qc����]���b�G�]�6la�|���9l�@h�
�N=�T8�Ά��Xs`n4s4�����Y��<�s�!��by ��
/}l�8s�t���������ꟼ��s���hW�ĲUs5,F��4���x 
N.S��g�߭ ��/��Ѭr���%F�َR9h���
�4�1��^&�h�rvz����
z3tio7���s�}��o��L�n�b^R�A�ύ��}Ej��}��d�_�^?b�����i���.[#j�ڲK5CCJǗ�d/�Č\%]\\^@�HI5���q�q��-�_8΅t�R�(3@h�f)v%�At��j�;�ff�I�}�,�K'Ng�sTW$�����&z����us��~t������O�Vp�[j�tH<��󱛛��_yr�%%��}==��MM_@�m;E��vvl�������t��	hk�_!w�-��l��'�QL)�	"L�R�Z���MܫTP�7�I�R��&@�hȲ�/s�(0��B�����n����������	200((R��������𰼩���O'��<<r�Ԇ�B��d�^}(o~XÙ�s$�tE�C'V���2с�6�#i��LC�	��T��
�� )��R]M'***��5@f|���4ʍ;�Y�r{y$��V'MwU���$]��#h���P��V,pyn(د�w	2�?Hߢ��q	�8��K!���M��Y�S�]ᘬ�dy��n28�ʲ��`2Nx�g��`����{�S��w�PQQ�>1!	�7�y�=	��'����#�q�_��L�L�@,���g�y��ns�~y�{�"/D�Ɖu9sĶ�(��G�1H�٤��V,g|�rŰ�>Wj��N����|N"����qEy�d�ve�w���8ǣr�P���|�[�$:��%�.2�:^��Ja�+Ǩ���OhiG���E��*(�22(��W�/}:��&� s�k=`rQwvrn���< ҹ<ۅ�ıeK���3��<�@��-�D�OP�����C�wu>��G���V�-V_�����j�}�N��33� :!Gj�#�?�/[���/{{{�y^.E�"F�EH)�ϻ/�^�1�4z֯��y�)8���"�h]<����DoR'N�Αp����Y�J���{yb�$��XRR���#y��8m�jh�JW����OD.��.L&�t�Ugr�i�#ț����:�r�_�v�lӏ�=��4�]��Y�?��vZ6�f���.�<� �ll?Á&�g��o�vC�}�����eQa�eoϧ���`�����غ��@@��y�^Ӯ \����V�F��9S�Ϟ~�'0���wH�p�	܅W��;522�D�
u������e���u�V\z��'8)���Թ=&��:5%/����/n𣥦!�%XT��x��*�ۙ��ƧME�x��$�"�;5����ki>o��:��������*�fڟU/�����t�����bnַ���e�8!A4�+�DX�
11K� bWr����&sf��$���#���H�~����YK[������O���VR�4O_����h#9��@z�#��B�]Pȡo�9�%��1ڵEq��o�^_H��DQـ�镌������y�(|�Ή�$n�4=��G���}![W�yG44K��'�H�0"ɔ��anv��h����*�I2������ܒW��� ��1+�b|��ݷ��o$���)�[O��%T�C��R��p����Po��B�����_=�T�#ݕ�x����]�T�M�����r�s���������H����V�c]_k0_�(��6��*���Ś2�o ���!^'��$���u%�ώ%�Yv6�h��������r��ݴ~�n �m��̫��*
WW��	6����9��N��C�O%�s-a�K�z�@�4�����W�=JB
L`��Rs�Q"����A�_�8�>c2Ȳ�4�"�����0��o���`:;��M��p;����[��LXJx]i��q^!GL)�Z�g/b؊����;'A[���F�La�bH���4�<�jY]���I'�V���߉o9���d�(�Ty;OeI���g����8k�l���̿�~��?�� ����b����_S����\��b�6؈gGfX )��r�gB^G_m��S'�2}�K �4����}�[�����'l� <�D͑B{D�?&Əe�'�V5�%��-A���:��ʅ��K���(D��Df�J���2ٞ-�D�5o F�������9?/�ٓ5��#�P� �!r9�-���ڣ��1X�I"T�I���[�2[b����0�l��U��Ɩn6N����S��F�U
�/p��?_@k�QMZ�kS,V��5k�đ����c���;U`���,(����T���Si�}����p=�o��!��Ox�u~����]y?�R���/�>D�UN�"v��Cb22���>%��z�(]`��Hg9��4$z����d���yiZ���v輆3�s�#�䜄����gXM&rkA�,0x��_��cR�9����Y��u�@��<�)��>���EB��c8n#Xde��� �4H���1���̐�eDe��K��8_�c��nҚ0��ʕҰю����W�;=��kX�с)�Ұ��`��,Sx�:�ƞ�'=�o:��o
����h�G��>��z�">_��^P���>B��_��N��'���?���o��Rt��o��j�Lë�L4�憒�Rry/ﭓY�%��\��u�.]����%�V_/\���ཤ��]_4�qMi
X)����B���
�W^�7]�,'���3o�I���Eݪ�l�CBp�ա�M��e�݌����Qz��=w��d���b@u�La�55!�o��FK������ip5\9J�� R��?�q�s�X���{"�F�h�Տ�~���i�Ǆc�}� 㪨����^U�"�O�	��|��yU5��4t��ce��M>�!l�R�� ҲM_@��kB|�ic)�lH	�M1�|�#��:q}���v��p�H�s�e��ߺT���BÍ���Œ@�%��Mai��p�J,��m�ِ3�W��ۓ�-��G�{�(fp��ͱ�M��cؐ_��`}q��.e�>�\��q�����q��.�ީ�) ��K�t����ˊ�oeH��Z�S���H�S�t�6d�Y��k���{1���&�_3�_���+~4��l9��o{,�s�-��a��+��W���yix��!/{���`��{8��yr��~����8,oED!��S/�v^n�8C���sz���%�_�Ѫ#�$6�l)����	��Z��,#�'�9�
�D��qσ�Q�^�7z���Ȝ�R|EE�T)���X=<P<��ӑ���]���rG�Cc�+s�!��¹�����(d
�)@�������R��Uj��RL��>�=M'\Nfs( 	��R/f�G���#�Z�e� �����g[2��H�����Lb�W�]9���o$5��3��qo,�zh4��8/�
��v���V�� �t&�Ư2�Ծ�wa 0Cʨ�x�^(C355�_�<��+���e_4�W��թ5k�����^����[�P�e5V��6Z=Q��\w�G��bd�ߔL�m��S�D���H�������}��)ޡ������W�R����R�N���I���(;Q��{������R�q3:�ۃ��+����yUɥ|� ��+\�g�������4Z'��o'`���uK���z��j�TU�5j�AТq1��f�L���EA��\�W�
|SA_t�I 8�BQ�$)�O���t(*��3��u��ᷥ����
˘�����s�[9q��iq_��>.���w�i�ݿ�FN5�,N;C�5��F$�ewe.=v����k��o��ܛO����Z�n2|z�q$\"�#�ʑ��5+�Eo��%7%{��t�i�q�a;�v����R����:�tI*>Ml���<��q�MݖF lt�Yȳ��h�����v���	K�%n���������K/6���Zh�������>�-i�E휟�5�NO�t��%�3�O������vt�tԏ��Uf��/2`uX��԰�0.xp��͖��2�Y��R7��t���Ł�Z�S����xM���L'vG��P��ox���#Q�N��,��ߍ|���)�t<�RX�A�Y���M���7��MZ|r�+����!����.?=@��Pf�UK�v�|Cb�!y����h���j�ꤏ.W��$�6��"�cï�T0�۳0|�����kȘ\�2�	T��(J��i�v����w�`���t�����<V���w	t��'�߬�vj��=v� ����>G����7�yh� ʸ��Sū�G���M�T_b�'F9h����Ȥd;-��V�!C�y�k�`�iew夛�2��`ʎD�����O���Կ�ZhP�Q�;XP�]�6��1�  ����8�h4-gմɍpl)趾��?��yC���7�h"�Qeۍ®������*"G��S��X�8�J	<2^Ù�G�8�s�S�]:廧xq�]���P�!��g����,U�5	��l��q �iU�l��z?�[��<���^�ql��3�Y��n�"�1�*�<�:t��
��eG���)����I:�5V]�%ù»4C3�]�+J�!�l�:IgD̙
kB]o��p-�ㆨ�C�ɟ��'��j�c3�q	�g�P�rEC5��h0�ق/���H}E>Dw^jaB�|�(�=4����G2+,=��S2IE��7b�2��y�sv�hu.
P�	��w}]�jh�K��2J�^W7�7|sC��>r���܆R$ ��év��#�&6�?@�(���p�iu���!�g��<s7����7�tɯI��N˛a�`'�+���"i�z��xXw�{[���OE��u�<g�kwOH�ώ(�:M���lV�Kr'[����[k��mdS!�c��L(�/V8o���q�9l�Vʥ֎H`@Y����ʺ˘&�I\ ���������(Cmp���Rv�o�7�r�Z�n7�i����4ު��)��\p�:��a�� X dU(Wd��`�IC\_�CS]�D5���P/
�0�е�S3���{�A�>$�뙕X~!_{���d���D��ȘjEc�%�ދ1R7��e'��k3���4����Qx�W�1���P�z�#s$��Kw\����4���!���g��+?����:�ܑ�7�[o���.{�3ȓ��7�� ��&�:��&h7�����)^�x�w)V,8�Ж�N��]�MKq�[���.������ߜ3;;���<�s�٥�xHVU�uj>�	��{z�C�UW��h���$���w�\�i�m�������:`5u���)���L��1�3�j���_��g*C���ݢ�l�V= �o���Jnj���`>OR�o�-)n	
j_��ޥ�r`���OS�]�Icd�e�+��Q��� � ��`�TJM�t�u,��Ȗs���YlOg���Da����(��#����r�M5�[v7,���M�_o�3�[�*��-���8���Z&Յ?x�vb�w�L0܆ ߼�B�����q�@nW��N�n�;d_�F+_l��/� ����D��ݲ��B�tZ�6s�I��7���I�H,��W=������0�Ҷ��D�=f����1-?��G�Ș����w�MJ��)u�� ��lH}:�/|�0Gr�4e��|k�U�I�Y�6��h�aC|�wB����� K�/]\� >��P�R���`M����4y}U�MC��6���Ns�<�տ7C�p��n/Gg�B2-�.������
��ُ(����#y�@�j�.�R�?'f��;i��&S����c^�l/��2Na�\���f���Z��u��CD�W��n��	G��Xe�߆U;b�1>oe�%7�&#�}&.���-i���]E@K#��PϤab�쥌�����pO�*��+0
�qX_��ܬ�9��,�i�l��a�M�gh���і�J��B�Ue���4_q���.N󅓈��;���c-��t �|B(����P??%姞����%:�p�����W��z��E*"$�x*��e8z���w3zZ5Lnk.f�h�t���H4��ݙ�kr�1W��Z���[��ȫ��i�����X�a���Uꀑ���N#x���|w�0w�ɹ��B{���M����ѐC�/�ʐ�� .�4 �����f!?Z\I��E������Y�lZ�A��U��J3�C1Ku)Z���kX�\(����;f{�Q�oM��(Z�P�-�6��b��F1I���M}�k�g�qvI^��(WPm��=)��jq�{C�uK��L6�/�cWEf�hq5~��hI�'=*�4A�2ǶsZ+#������QD���G������?�i�U���g^���8�֞�����"�= y><���Ξ@����{�;��];ЇY��i�Vu�#?�\�.����6�T*��L���+����1Q�W��m�v���4&�)�a���D8|��c?�t���?�El�d5�**H����A�|^���ğ'n���]�[��#�K&�Y��	��ٕ�6f���j�]*U�]���������b���u�_����$�k�a*c�F�\7��7_ֱ�����O>����T�����	�Έ�l�;�Ph=x�o8�����/�⏙������b�A��9uJE����$����eY��4��7�w/,M��BC����<;	 yjYF��[.�-�����0�*�����Oۇϛ ߾�4�|�ӛ��T��G��U��O���M��E�i���M�~@?f��4���N1�MQr S�v�ڬC�r����x0��Rq���gRO� ��ׄ����HP~T����=�����eH��I:bs] ���i^��V��T;��ϻ�*��}(5M%w�]�aX[�5�n�����S�k�n|�)NJ��%�bʀ����/�"���7�$z����đ�Rz��a	Ξ��.J�­J F������Y��]�-$=Ν�����:΋�ɷ�������6�b���O΂Yi�9��S��<����`"Y�^1��-�T7^�Q�/7?Z�}�C&���^Č�3|�����BQzѻ-!��'ا��G����l�$
�(6sH �
��[g6�s����ɡ��'笙��Z��M�%+/�5�(.��	� �Z4�����x�31�F8B\^�?���DDDj��?�	
~OL�{w}������&���E#�K`eeeqwu�wo7[?Ń��Cg��3b���N�o��u����9*�M����]��Cu�DX���XQ9�����;)�d4M*�d��JD�����$�\�r����3��:8`��̋�Beł$ �$y-f���L!��W�Gҁ7Х6��ҹ7�l��!�W�+����e�:�p)�����y	��|����2@peH&ǧ.�����U����Q��?W�?4��NUL���=�熭�r��W9>���[�֖b��;lu�\��f\5>�H<���_6���\��O.~�}]�'�'�����M�a��Y��tG����K<�%��M�v��o����bCE�Ϧ���	�����B��s�o}�"l,b���!HW��Б<:� �ǻS|�&RRRJJ������J�]��冤$���7��}GV�nq�̻��F�C��1�"�2ŷuϳ#Q@�}��H�rwN.�F�f�	d��%�i�c��A��] ��~�	&9�I��t�)g�Z9/��`���+��W�W�l��å��E�4^�����2/3��h�RG�K�j�\2��͞	��nY���xsFd�Ǥ�Ȣ���$���>�m4��������c������M:^�.,�]<�Uw�'��૫'~�R?�Lh�b;��Kf%q�S�����?Z�[��}-��|o��������fn�~R��������e���A0S��P��.׫�u�0�/y|���]�V��7�	e�CɏX�B�/�p"����&��^�ä��s)$��aQOg8y�X_��8�tfl}�+�V��'��?S@�
�-�1Y�:/ �Z���M�q3���yr��m	J�0L���D]Gٱ��?�l���WK��������~6�T�HD�6���8��"'�����^��*vR�En�6p?��e�������_a�A��3͝�]<�t�'�c��w�LNk�ݙdB���gm���:��;U��__����>s�<���r۽Ei�e}RfQ���X�ܧ�A��l�K'2dO�	�� �Mp}��d��w��X��*��j�\��nol���UXUX�¤T�epP��c��������<�����27ǋ�j��֊��n$X�L8WϹ���Ԭ�w�>
��7݀W���BU��f���&)ا����4Pq��������G����7Ç�1�@��6(��+���*#����p2�	G������R��ͩ(��"��I?�l��}8p��c��B�%[��ɕSΕ݌�F-�Fȉ�s�Ś�Y�Ǵr����"�S��l��R�k��K�5�D��ո���Mm0)�^��6E��߿
o�ؐ����Jy.����v�e�˨��8OOO�c�P}WG-�pP��J�}�Ù#;��Eჱ�!��sb8�ծ�-c��؜w�k��O�/P~Et�;k�j<A�w$�t�/&�V%�*�2Aw?�f� �)�K}ǣW`�W�0���0�p�ծ���1�"[�~�9JUU��ѝ����6��JcV�β���s�8����BgoB�����<�X^F�J�F�i �p�Pӎ�hb"�q�~�~ :[�n����Mz�ҟ��=p���蟢`��������>����7l(d=F�=3UWo���(H�~��o�;���l�7�j����^��8��vlFA����t)J���ꠘ\%�u*"'�*?:1���@���7{L�k��D8�(��|]yydTK��ꇗ7�Ǯg*߃i���n�쨼�X��
���zZ**1��7�c�y�?3d���F_m��w����8O����ز�4$(���f���)|�c�9�*�4�V%�ߐ��舆\���PhZM�tnnn-Sӷob��6�=���;;s9H��{������������1n�k�HsP���,�L��Wx]�Cz��!��t��Š�	���
�/)�hzx&�(�����/��YYY�#J_�+��?�!��÷/��P�nz�
Io{\��{p���R��Wh����-�C�4�7a�/N��f�m]�����M�<������~`Ց 
9�?�^,���� 
#��Z�g�M�F��=�Cb)�!{e����� ��H�K�1�a�����:y�t|Vir�'0$P"�!��	�E���!�DX[%�Qm��#]���l���o�\��	�Ì��p��80��M�<�l�,/OS�QT�~���grk�(R携$�'�7̠x�X�R�W��2��� w(�v��T��ݺY9��X�&�;^VJ����xʝ�Z�: �մ�!�U!j���>
@b�'�E�jp/�u#Z��v��<6�$��^T�Q�vG;��W���E�C�@ �K)��8��i��х�f6���3�����J#c��{�n���HA�ór���)9�U1X�h�G�}��F3[�,M�aIY2���[ng���r�nt�)�R\�g�P]S�b8�H���"��Y�'`,U��RG ���`�z�v�[m1����
��x*�6D�#-��[�X*^����_e
�����{�E2 H$N��=(B�^�z�~B㯧�'Nh>�ǲ�1���o�
Dr[�1�2���}�:?b�5{����1y�j���ВT!=����m�Nڹ�o9��NX�wr��C�ɟ5�K٭h�+X�5�e�=��G�.j,�~D�%2�m]��<Pu�N�@ʿ�?3�:�P TxNayZt[��<�פ�`.֪�q���y��Ɉ�Zu�<&�����Ub�0 ��;��ՙW�C=5���6~od~�*¿�-�����әB7{�r#�5|��}0��/�-��ѥW܄�t��;��=Q�f�\�K�f�����S�i.�D>��LM�T0Q�f!��5�)�d���;y�.�-`�jX�_Y��9�wN"��\m�ұ�\�����ʽuWѾ�p;u�]�L�i���	kz��+$5���B� 5b��u�Pa1�K/1"/D� �2�������çTo���vOxNa���R��D�e����z�ng^�T�����W1����M1�E��#EluD!��y["l��X��2��� �3S窼Y$����r)�E���yHC�������<�N��ޖ�XͽXDZ���(���/]�����4�|�ӹ���}������ �<���1Yx�P)Vg9��گ�-�V������"Ү�~f.掊�e�������?��� Af�p��pi�ᔒ|�ک���Syz��`��s��Yl�P�����ʶ�:����9�����a�H8d��gϗͥl�oG��� {�]�$%�vJ��l�FE��fl�]{�&�PM�k�1'm߸W�Rt�|�rw9e��Z�'�B���[���	���xRc� *2m�8���v��dRb��fpȣ�����f���ʙ�|TH?̑�Y|��@��I���+ݤI�}������f&��hkhbh��p�?p 6���yH�b��մ>Cї�,er��V���d���z�[����2�X)N������r��I�vBRI���^�K�lBhf����3���n���"��wܱm6�o)���f��P/�I���7�Zl�a�E\3 ��rs�&��T�%�/�X�S��:�'����onˋz<�i5�Y����PM��q(����\2���9��cϹ��{�����H�(�4zȻ��?M}��[�e���������ƴq�t��vu~/���CmR�w���s����M7����5�yo�g��Ŷ��1l���*y�$=�$���l�U�PY�Ey����W���rĔ�q��kj0/.'������:b~[�%V9�B�7���6G�-�r$�N�Z�z{�b�t��սj�,�j��6�{ ����q�l#�-i�G��3|�-L��c�Ꮢ�4� ����9�Cs���>�_�U|o��T�_�F�^q��Lz�h�Q3>_�\/�ɽ��WX�1�}U�	m���w�Am09ɬZ+H���ES �s�P�F��?��`:�#~o�߬%�~����6�>N�@�3Z��xWӈ�6�lՅ�5E��H�Ġ.�>�T%�-Y��3�9�R�������XN3 ����0j�E�/|u�8|bf9ī���x�p��]V:��c2_��9���w
bކ>g"�P�g�H�zX��������P�/]���WH. JZq0;l��5�ReH���&�&��ݗ��}O#c�ͺ�����E�4�����O�f��I��dU3��Q��Y�����5�?��`�_���yv�)Ł���oA$i��0w�����w@B��A�p.�;hj�s�vl�M:���]��wB���sL_��b8��~� �|b.�W�z �~�R�y��L4�2�W��fp�t�`!�J>�����h�[,����7�[�	�<EiG�6a%7�:FJ5���r�=s��_g�o�T{[x���'��Q���qȝB&�o�Ų���`��z/�8��;=ץ��L����i�0n��M�{k��Ա`�E��j>r�7�	�_`�ÚN�\��q�b<hm�����O�E=����v�N�B�d����ڐs�e�Q�[aʴE�DB���E����5��<�8jSy�k�b~ҵ`�Ԝ��$/�?V@X;��W�s
��}��� $�O�Ց���v�m����U�biz[-U���;�&�����:[tw��C��l�����'j��Ix�h�+�X�J�1�2уP[�fxmX��Gw��o�0B�ozn��D[/B�Cl�+G��j	�5�pl��^��������j���h��폗�����g؎7aY�D�,��7T���I�����S9�,�8�l�����E���o��9XN1.{�}�z�E�	�)r�,���ѫ�%3��S�R=�	��?�~�܎���B��L�\l҉��;��;'�sr�?x.N��,��>(��{��E�l-�%�)����^��O�Ǧ��d;�_�V�/��!�7�-��R�@}�]�{�}	��/�]yW�xH���N���{އ����(����������
�ɮ�8�j�����*fQ�y�������I�>��L�./1m�6�B��٧��I��,3mu�J�tޜ�鯫�nn�vqa�ǵ�i�a��1�kH�uWȊ�3nb��ȫ#Vo,u�oRan|�y��
��[#��D����$i�u iE��5&]t1��U�y4��<)42����~�//����W]���>u���H,����D.���$@�K��E��C�*�U��^��k�{��"��]��K�<^iњ3��_[��u %�l�<������������g���a�
e^�������x.���V�(p1�N�4Ê-uS��f���/�����}��-<>"�{]��.u�ܶ��̘����-����,dPN��0r0b�Dc�.��Z���!!�=�3�k����᫺@�F���鼰�׌d�e?:W����p�=�>U	ݮ��|UZ����S�r#�s�T4P�k�ltȸ���S����NWP�ݝ�"\���<�\	����T:�O3Q)Z���g 3��g���5� �F����0q#�����b�B�O�{=�嵐����M�z�F_���/�����I��^{Y��q�/�Z���������J~('���R���Sdp���׾J��q�~*O�0�Od�U�4۩G6^yi���5�c�*���
om�v��&��~iZ��Eߪ�q�$��_@����J�[7�����m�*��1��!㏦�=
L�X�kҡ���i�\��A!eˢ	��D�~ ������ �gH%�Yժ��,~~��Bs��08��<Ь�ڭ���2�"��Ǯ����[���mE��{kr�3U^K/�'�����]3�G�3❳T�͡��f�v=?�J��m���H4�z���)R�تq_3�߸�RB���ڰ�����A��m����<$�v��,����	zt�qzd���&�e���O{���%���0%��M�Ⱥ�ՠDg�-(�8fI�7Kܺ'I�x`.�?���li{�H��r3�*�Z8�cC�/�
���F��7�v�s�g�H�C���ǕT-3������6����r����8�s�lז���h0��Iv����۷��w�V�-h��X4l�e���mG^�h9Y!�,��O�}��>NʲA\s�Xg��6g�
��w�c�,NԿc��X����� ��E��8Cr�v��ւ�'m��h��3�f��,0�l�L�]��#Vv��M�A<��e�Z����ؐ��˫T|8
�5b'٬��J�7S��e��o!Օ\�t[�0�+�јed����şE]J�Tq(3�@���@�ECS�h	�C*O�tGD ���� �{	Q_:�G��_�^5� ��a#doA�!���,�f���+>/A�UE�#�
Z��,#������ �1��K��M�Q+��Q.As|/�%�R�J#s�WoC�H^#A�������'�"PQ���I��p"� ��no��r����Ă�;%�/���,�E�gxR1�/���1w�i�����[��%���_�{�yKWK��?N�x?e��~)X@��x��[~��.仳U�/k� h��ee����D��w�'u�� $ Y��p���	@*�)��[8֕��2�Z6\E�g��bL$3���x��o�3F ~��%AiT��r�)*#cx�<D}� H���Ӫ���dS F@C�j��?Ic5�8&@z���'�a�&˟��ED*��Psgb��K�P3� �4:'��l8����Ϲ!g���/��"��An��3�����?K{��l?0��̋��z�tX#��A���O����Z5���	E?��11�鸝Ey��`��g1:��6�0ג3ڝ�^T�Tu�h��Y���Hw�!|�eZ*�8�������Q���������C�0�6ʭ;�H��H�j�*@z��>�H�DnO�ʣ���{��$��N/`�8]�%�׮��l�w/2A��
fŀ� 9k��+�vp�_#T�� /9o�~IH`=�zc��yM���Q�ğ�Q�|�<���/O�s�FH��i�0��R�F���V�W�("���"����R ��O�-��}��V��OZ`�?�����R~'"��4��܆1��߿v�+"��5[(���y��H��pٍZ\6�[��U�ȜcQG�0</!�x�	���2��p���Jf��}O�3�FG�U;k��b������Yl��	�?�~6ϯy���	���7g�l�9J]n'Q����x���_�k>��K$?�y���;^v�n�{ɑ�J���峲%//C�����V�N\�L}�����ۚ-����[,�W�������~��K�-��F�y"0�A�';��!�VU�H:Q[�O�k�SWV���DgA��
�y����s8��߉!��m�Pf�<��M���}2������a������So��%URE��a9{K��/~٠_V���o�E-&�?�2�a�{fU<m�[fh�溛"wC���*Z|�Q�m?r�\M��c/Sǰ8�]
�浺�ɷ��9}�*�L���#v���Z�z5���<45G97G=��`�w����C� 6��}_k�s�?�b��m޲�����K�a7�Ca�f�{_X�(�u�Yo���a�I�;�x����Wa��a2�7e�� �c�!0�����������s0t�V�Xr1�)��ÄA��1��7Y��I�H8mo��ǒ��L[������u�Z?`yܳA.�C�p�����^:9�PY��6̤��?z�M�k���1�eB�	�P&��P�8Y�<XL�m��\�_�B)n0c,��NŰ�u�}a~���,�X����!>fCc���L���]K��f��'���aRVNXp����v�W��թ����2}��a�u��P���j(���o�U�f�8�9���$��-��*�)�_���ヶ�ﺃ�	[�q}����Z����Ѣϸ.�S�^�kJ>mNM�v�Hv����n�j���Qj-��7��<TR��i��@�]��a-�W/��[�	�5�4�+��=��DΛͺ����bQ7
�.PD�8�rƪIFT!���6]�}-.���M7)i�s[o�}<���ü���D$����	m�6����@�cmQ��q���u��%�GG#
��gQ�j���[�S��Q�d�Gpo��~sn�_3�l�� �=��ʣ��;8Z��+&}��g$��SXq���@��������]k�Vz�$���U�;�)&P��$H�<��F9���`��x���$R�4(�c{�p(`!�4R( 1�ǖ�}6q�?�D���2."���MA+��62q/�<��fV���(�2g���& ��D!�ro^�e��xV_�t	!��8S��qWqkz�EB��D����F�K!{�L�U�]���GUt��z�ߥ�1���c��C���ȫ���t��0��u��=&|D4$���ǚ�(6p~�|}?;�1d浚�x��i����1&.���v�06@��Z:����
���/�ƣ��8t��@(�Y���g���O�a�Tt�`�W�G�%S4q�Q�.��5���L��A�`X���_X�=���еq��~�L+ִCgX��5aV#>�sFG����>`�֔����
4�b��"�·AQ�WcB��ݜ�E��s��Da-H�o���w�cT�2^�d^��(��<���lòj>T����#P�%���+#q���A9�9o*K��A�V��RK�>����\Ca%�����k�j��f+�#��m[�w2�x����J�$�P�j@fݾ��,&�c��d�K�T��қ�y�M��_PnN�l/�E�uu�o�n5��g��1���m�`pΏOE�� e����r�x�u��L'�G����}�X��'Z���Y�hcm[�Β�5P��E��Q�pw]�E�E'c܋e��;ЊՊF��g�L�6*f�W�3Kh=��jY�J�O>�����G%��kӣ'�+|����T}m_j;2#��O?J���ߐ<�:9}mZ�;Md7�OB=6�>��m����Tp.N���7|AU�J1]B
(���5�P�Bk���kGeɟvN2M��R���M|�Q��)�9�g݈��.�o[؃iz�wl�ar���_̑sCߥ�����;��|�D����:K�����"4�
v�}as��@��6��{L=}1!(����$I����G�Ja���m� !��+3(AD@&���I;�k���{TtM�>$���P�=lB�]���S�U�7��=�k�"�.��� ��g�+�1'��������&ν0�Ԇ��Ə�����Yc��BG�V|J�M��&?ʥ!�z7=&N�&�~�#@�=<�ɳH^>c���j~4Z���X�e��Xo�3���ڼ��p���S	=�����6Ɔ��z=4�^�!��;t03�k7�V#�0��&�/����)���X�+vB>+�z�w�Pm&�y�J���x��.�QdW���J���6�FPR�h T���&���j�U���N��O{��YR���9c��Q��nExV ����~���`�S3p��		>{\b6���7��F�5�dk�O�O�\~�QIA��+@p�5Ɛ����,�b��G�t��ؙ>�GW��������}%���<�]���^G���^%�8�]{dH���#ڧ:a�N��UFqb��\\u��a��%��#��L���C��)ST�\�F�W�]��Sp��g�M�= I�	�P��;?��*�7:����W�+~׾xa�a&��?�-�Jx�X�$��� %/�0�F��o��?_��<rZ�$��}����:�I$ADĊO������Yq(�����0��^]w�L#(wv�t�rѷ%�ٴ'YG��s����ϻ;���_A欞,s�7��ln�W4�w��&��S#�/��@ǌ�Ir��_�d���~巙�W�a�&�r�f��^�xF����$*�*��{֕&�ɥo���$��	�l-�!�/�`Ҝ[�Y(���IS����&-�������O�l��Ou��'v�÷��c���j ����(��#����y襜�dփNPFr�Bu�~�,��"����_�=��?+͇�M�*��!���6� �)1酶�@����[0�w����V�:�L����͍���������x	��*�8��w3W���w#�*�:���s�W1^��^��k��`�X�I�����g!EO�J����Z_�KJNP?��?�:�>`�߇� ����"�IƷ����Xe)��h�����ev�~M����}��Ԝ����y+�&�HG�jE�^�nH]y�,Jd��� �����c��~�t�@@��̇j��e_�<���yD�����}t�֑�)�<��P'F�$����)�Ǟ9��z����OxJ����|+�G��(5$?dj��W�8�V .e���3#����)��K*}�f�~G %�;tRu�AW#S�n�;k��v��%��.���%GsRξ�s��	qMi�U�@��l�G�?���R��%�۲���мW��:��.Ţ�?:��j�r��ӳ�����ϲ ���˴¯Ǽ�m۾�*A9���$�@���4� �(Ԥ���}���vB�zBh�&������T@�p/��ډ�R�ק��T4׮��~�;�'�]�9��e-��A�T��5�WW�����sA��r��x�8����s AE3��b��<���2�Z*�����퍒R�x���oz�, ��<��̺���5�;2���Y�U������ ���C���4Tr������7���u���D���W�ªҊ
��sݸ[߹:��VNA܁�}��`���E�~B{=��ob4�LC���3����nnfCk�J��g4룞Y���׫o��]w'qo�O��_���؃�.ݚ8�ߥ�����\}O�&
��@�"ϙ%y�H,Ю}J���{�y��_��Z�9 �A	���}�
A��<j����0z��cM�{��7�Zf���ZI�_���Ԃ����IE@BF��������A��hw�#G��c�_{��E�e/�}k������g%�4��&��Aru��	�\��p���S�bs���&p��/����d�Vp�{W�'�'�� J{�Ӳ%�����KJ��Y�C�ȓ�-ׯ�|!	�8XX�7�]��xh�U����乤w8Kt3�<�~jx��Vx۫��޷0��`bbR�� Y,�Z?Ӑ�(����b:u�A/+3�"佹�Z-�����$�)6�n�$�&�T��}�e��[�m��y��������%��$�i;�,�3��I\HH���v|tE�rXjm�E^~��4;k0�,��t8$.(�||��R[^�����ˁ2�'q�H�KAwo{�9~dEi-p${�\��$��cdnn��=�6�
���CCQJ��$ֿ�f.�>]=^�}��xs>)�Xk�0�#���0<n�·/�G�xl��WUW����͆�Xf���ڈ�9$p�u/W�*�ܙ���#{5~r9����،ߌ�10��v�B�Ҩ?e��U3��Zt�����r����z�i���/8��I�!?���o� Lt��%҆ml|H=�IT�i����m���;��L��#Z�QW��㛿�n!,B�$��y�9��J/�#q�ю:.�}����1\;�S� w��+x� 2���O=C��=N����:����Z�����(�|�٢6J��`��P70��'X��fg��3}k�2Vg��D�qr%����"���s�ԶE4�Mj����+�/��q$W�||��������L�,���?i�ҽ��҇K�#��0��^x��*w5��'���c��oR�8M�G�����ut6<�F�ٿ ���P|R��oVu�=hv{ItRVuF��	�c�^��B�/���LMiO��x��~$X���+����e<�C�'o�����]}�WF��6��]>@�O�D^�IL.����U�W{�(��Q���.ͮ����D��|�"�Z��}��|r�>����tfp5�oΟ�����m�D"P����'h�fzlBB��"�6O^��^<�'<��m7�5�*�2;��V�Z/㥚��i=A4]��U�y�C�c����hD�D�7l�	W|����N_�
g�]WY�6���M���z=� ���%���+�%��V�䃔f���r����q�[�������������n�`e��Ȅ3�,������U�A���M�B��b�w��|\���M��G<�h���r���!�o2!bQD�]�� �qo1���.f��a:}M���SPZh�s�,�2� �:���ǈ���	:����Fɼޞn��&m^�|��5|�I�,�Ϣ���R��O��
_"�~��Di*�i��)N�R��F .��8b�K4�+zT�'zTcv{x�F!�"��9"�]#>�^ՙ�Nss������RCsR���1�qr���rZ\���3Y���3�A�UFI$�4�6=�Zj��`<ǋ['A�Y�rH����>��Q�&d1���%�1�l���2D��q����oN�|Wri��A�%����m���iԜ�zs���7ʎ�����ǯ��<q؛���~��'w��5]�����@��� .�_���)W����UWp�U��#�H������/��QN9$�|^��Xץ9�TP�[ ����z�?�����4��m͝R��1~�.ӡG��U�~G��׋�Z~K�2��G`��C�YQ�ٲ���w��ׂ���Sr�e��/Esz��4.� '���!�k�
H��~�㟹]D�ls���T}>��H���g\z˱Y��`򛟉��/-�.���$�DgS'ފKxo6ߣ!I99p:b�����/Z`�hI	G��#
G�7,&9
�����> ��l��,ƥj*\��n��Ũ%j�=�E�:Z�]���B��Mi�R���~�q���4���Z�w�\y���P�${��ޥ��Xw��*P6����P@`�"��������G�?EQ��j���cr����@����E@R�Q"=�4�Zg�,���Ro`��i�=�ΰQۈw�^y�P����0:�z���VᤨQ��k��°qO=o�/�]����lo^��'�0jL��?��X����/��C�jӌ�z�����q1C��%y����JCĘ�e;�y�3�B�n'YQ Uk����|���_�dC02[?O�̀��ݎ뿞`��#��6��-W�8��]�� �A��i{�����L�u׌��������Ű�9t�g�.[����S%��7���sx11���  ڒ�Z�6�����kp|��P�H�"ȅ�����6jA|���c�a����O_��w2ˣ�T��K�+��'����[\ }��P��pf��;��z�?o���L����g�W�K����7LD��10�ͮxv��O����Dn�+�+�V�d��e��ߞ����K�()��Լ�"�;*6�U�#J��/�[���bIE�
�#�,�5�z��%h{9�\���fÌ*�WE��ï�#[�T��\�`�����x�/�y���q'��o_�^�c�u &�T�w�6H4)��n�>�ڎ�A��Hs��Ʃ����Ϳ+a�z~��c�E��\�@��+cZ��eM�n��5c�棉ay@�?M�&@=�]$����iŦ�Վp�=�/��F�',�xo���\5��K�����cL�Gi�waω�mGϳ�1���6���&�K�?G�~��	����͢zjN��p)%3Y?�����W���GP�^͛G�|��\!��DvP��`�#�~��$pY���C�7PVu��*��cv���=�<��pP�_��1L��Qp�0�u�cx_qE�m1���ߝ�"&5�� �:|�g�Vm�4b}%����ƪ�QZ��0���b��Z��<�R\�������[}���O�m;��(AY-}��a����33����?�SS�r��l7��>�
��p�g�ggZ���:}�D@h\�|
Z��3}*���~	aa�a3&D}Zuoj��e���;������[��s7� ��s����k�����3��q�� �J����,���qPQ�W�C�*~Y�#�9�hf*�p�/菴����|�M�ĥ-���P^����E]>�/˝B1:h�t}�O�_��_�&����X�2�HZ�����ʳ �^vw|�k(� 4��E�܂��C��Ό�0"���NuG�f��z��<y�m���`�>�OkS����DR̗�?��RƳ�J4g��R�R��`�I��F�a��9�<u�(KBI3�.w�����^�
#��.�o��$�;|�R)g���Tm��l�QO�5kŨ��j�l)j�R{���+5��h�VT;v��֎��*b�W��;�=���s����s?���������k�`���������������(�J�Q6gl��_�O��.�^��skJq�Ht!XXI�A�~B��.�o\p8_it6,�C�>�|Ěrߴno;3�O���(��s��-������'�Pc�]eϭ�6��<xFN[�l�^�JAN��B���T�3`<�����Ѓ|2k�����\2���i8��igkZ��)n�����_k0+������.iF���-������ %b�����3$H���~�4�'*E3�bP�T4/��oy�7���'Qi�C�`���DU���:zK��,)^ʷ a��5�69)m����J����([/���󭣀��d�,]�\�[J�-X�g�魬R�爭,1��0�n>���pTυ�o@�d{�!��߽��,L�v��<h%��-1���/�hY�>�KGI�Z�1[e;���1,e����$7�(;�,.�q���F�d��3��IL�)y�N��`��8^gB���LV%��s;9�e����7���N!n��y�wk�s����\_��������;qR����P11��f�b������k} +(߳%2������2����"�,4�r��H䐋��:�$i%�_b���#�HZtoR��9o�Ҵ\K/�jܰ��Ⱦ}_*z���N'�b�����9@3b�!�Y�3��%�(��3+9���i�_��2o:�j	M�8��э����I�קQb�_u�Ѣ�p��I:]�����/���ɡ�qD�97�m�!o�f>*���ޅ�؎�rh��v~T�E�[U�qU'_�\�b|ٯF����ā�z�|R�t@I.��2��!����%ފ��@��j�h�_���;�9��:�K�%H�� |�-0��� ������Iɽ�ި���<�G^����6�i6%��"��v`����4���puM�w%>�������]��Y���؃�9��ң=��O�w��INob1Z§w �jP�e�3����A	��3�w�3���&ƨ��QGR��WϿ�mZGNa���ߪY]Z��N)�_ʇ:	2ᰡ�pr� �(�9P�(4ʲC�ԏW+����,����T�˂W������g�щ��q���n�s�B*�n ��MU'�����KP֧��,�4�7����:�A3��Ru=�$���Q�����p}"P"�q��B#��������0�ɶ��w��yQ}�f ��ը��!=�
(�A�h��]�t��X�+:�g�fa[��[�Q�u�<e��~�K�>�׵��������M:Xy�-�}���{��!�_v�߽�M�G.�+�Q����<dѭ�l�WŷJ�ȃ0a���������uE��[Q)�1�>��L
@���GPcw�1f�]���h���7/jUES�S�)�-���'�tq����Ef������"�r B��'��{���.�6@�g���,�@��Ʃ�MlU9�U.S?��ua1��ʇ���G��sLX 
:��=����1�<�[��_"���&�:���ӌͪ���\���A=�b�C���7%���"�:ܔ�,]��'�K�ݎ���GKT~h�14�'J�VN�2��d�3�	^�rP������;�L�dP�p�)&Dyo�J�8�ĥ�1,��#�L��\>�^{ы�zg^қ!�"4�o�
'!�%�'�@K;'�˅����y����i���};)��3�^�_�� -����|��u�}�d��T[/~@��f�8��X`�j3�!dpAe�sqѸ����\��-l��
��8��oo-�aB���~v6k�8T���v�i� .�n���Y�e6K0���0��KF���a�F{�i��[�2�h1��X���{͛�4����ד�����i�b���1l�^�4�: `&Ȏ�7͟��Z
��ٷi��\����u��)2^C,�@3� ��ev-:�Rwb�BҦƛ�a�<lVx~�(��!y0��������@6"<n��������'#)-��cO�f3�3�����]�loC8u2B��������K���-8I&����7�kx�Ǆ��� �F��Ae��:�s�T���3E���[��%m���M���i��{^�KM�yIC����|?�Bɉ�Y�d)�b��].qt�'�m.�[_��'0/�!a�2X�c'1����w/���ё̟�`���wl(���A��^����薕�^�2���(��B=�P7��c�s���ZP���?l���ƾ/e��iU��2Lj��,���]pD�F���ԊM���` kY�g��5��'~ܸAx�5���jG�ڀ�*�3�VzD�{�a�ʜ>��7%S�J�F�S����o�Xv����K�IHA����#q��wb� �v�6j��9<�(�c�����!�+�R�˯�xwL�j�"�Vu=U�Zi�/�\��^��XQ�R5�nf�=�3��_��7��ܲi�ukg��}и�s5g	��h����?ɮЏ<�O�Ľ�^ %�R��.(����\�`.�0Ր/d��5Z
."��ۻ�tmd0�Ll�MJ��t�:�+Z|X&����.#��P۲�b7"Q �?��:�B�cv��Ja7���T;r��m� N�'OV�$ı��F\�>,SF��T��!���ۺJ�a��S�@�ʔY?����ۂ��N4R�I݆��[�x]�M8?LN�'�߰����^25>��(>;�����쇏�wzZ2" ɩ�ʲƗ��^�)��#��3��۾2�Ɛq(�IW?9	H�!��xÁr�-�O�b0��oL
G"�rX�o{F禵��B�6�b��ve�`�0i�<�_�!.A�?o���xJ)�H���SكPg��>8�ƶ���ɿ:� +^U����ɬ�\�F��9��2D�g�������,)j� T{��|~��,��R�ff���Zq�X��ȇ���;�$�W�T�z�b?®3��.-~�V%�R�5A�Z<��u�?�[��԰H93r���g�/(���P�0�e���@k��I��	���VN�[���X���IqY9,T��+W�|���P�BM��`%.��Hl���8><W»R�7�k�6q�r&5���n.�M���?ҩ�w�Z�|��[fz]�ֲ^����(Pː���e60��`@�u�U/��'гR'b�\���C-���oDU0~��(QZ6$�#������7���]�Pkt�g��o��`0t�a5}�V���dU���Y�s������8��r	]ѥڒ�1~�*�����a�yiw����	)�u��,��[!"��^,1�t�\W(�-RM�Ҽo.Ƃ�l>p^�\��ؙ��
R��<�!���D�������*1(!��7����,�b:w��b|� ^O̼ٶ��)6)��y���lG�)�b_���sv�	�n�g��cʥS6Ĳxf
�qO�o
`�֖r���t�ۆP��)Gˇ#��ٗn��.( Ȕ��9�_B�G6{����`����u�*���n����/�Qy+P���AVfg[2��-s�K1���9^\�ڮ<�����ѫ,�P P���>1
�fB������{��ݢ��@��;�!O k�v}�Ģ_aI\w�ɯ�� �y��GCҔ���s��r�@�=�\}��y���g�w�ͻ�m8^&[k˵��+�~��k2��3ͻ�=�y&ϞpYVv��&ό�i>�#���� ���C���Nb��w^�����}�k�xl�Q��E[���<�<�@JC��5�#5�Gə��pwYއ]|J��L��eڸ<ӑ�nE�ꐫ����g7�ht�=���g��h��߶��b��pJ�fH[}!��1b���4O��DՋ8L�J�6[N+���*��嘮?hPn�BxF�$�ĸT���AL��u��Ե�x�(���S���NI�,����a��1�5?al��T6����=wp�zIDi֥�����MHd��W����A}a`k��f�}���w�"}my�G�r^ݑ�ƪ���N�V�0v5n`0Ť��k�Y�h���/��ut��.�~7ӌ�j�6�����J*��U����!X�6�="��d�Ȝ��`�]������3�Ȣº3�g$�}L���Bo��}�e8r����|2�V
���H�{�x�#X�7�����C���K��3{�;� D����j��C۔-F�N��1fg�b���P�V^������H��t��� %K����t��<�ZLeG��C�:�Fx�%q��=ip{�8�{�P������^��d�q^*�G�+z&sI��W����▷^ ����n�!gb\%FY�U���!�C��������A������\���Yk����^��!	>�X7y����>�XrO ��S��9\���>g�i*�{�i����3SMq��u��]�V$hE��5�Q�Ϊj~�5�2�Gb\��O����V�D&8�^؞N�!=��$�ߊ⧬�W�Vd�ܭe�W���ۚ�40R�E�(��:�˚6;�(j-�(�|�������m���If�T�GF��2���y;ߐګ���S�hJ���0%�=����@�����twl�pX�I�+h"���(�ߥ|m���A��>�q�j~�/���u��%�`�u͹q���9�A m�(s��ux]��Df@T���&�	O�����P�:q�ʂ�N��}uu��+���~�8ж�B֌�{ym��@|k��p?	�n+hD����=9W����̌�2/��߾�s���������[� �3
NJ�P�:L>�>� (6�=4����ƕ�Fa��ܮ�D��$�T���H�,��0
T�?�����U��c�<��7�ml�Xy+9Ѻ��1��`��m�qќ��Aj�BIԇ�rh�)S7oW��i}�싑E8L<7��
q���aF �Uʕv���F��l�Gw�����֫��
����
b���8�խ�E���� y�6��r�l�]�6�JC�[�yD�v�2�<�!})΂�>�$Hȿ����ëTK�� }��פ	�9�-��|��2�Ps��x����m�7h�R�)�����P\t�Q�!b�8��_�3�C]�'��D^i�}bA�D�j�tH������"@w3;�Ϗ��u�|Gx[�Q��@�uQc�X�I#zٽY�����j\v����B9�@�/#3�JD,�)���B6b(��k�P���L�ҙx %�*2���6*�2h"ӰQS����C��)�#��7}#3s�ǞkJ�]��E٬�\L�9���sd&GC�� �;�M��"&\}����Y6Ms�=߯z���/嬕����������f �����س�S0�s��\�>��'��v� ��?��l���+��~��t���N�����2E��Z��\�k�=�`��/��'��)�/�v1#ĕ�;L���F�g��<����u�>'��'��?�l�k��*��~��bEa9�ϴ|�7�xb�\�-�HOh�����r�I�(����9Q�i�!�A�Ԗ*�K͛|�nn��t����-G����j�4ǧօ59V4��%B9��tT����x�\`Eʿ(��.�?/�:%�lĎ����GJ��vnn|8ʮ�}�]��M��ۯz�¤�k������'����Nki`^���w�Q������B�JE;[���D0Iο.��g�m�y�~%z�����U�z*{�F$�*��~�)�����&�Y����Vd�sh����b��售U�2,8���Ϡ%��g�g]>�'�(����x=w_����֒�`�L���V�����X��9��_{��:S�f���P�4�U}��0�(;�*.��~�sZ;��Ī�ο�u�i�8�՘��,GVT��eE�����o�Q��o��!ehb̪�8
�ڒx�n��r��G�h����v�q�q��ϩ��: "�ʓ�����X�j��Z�*Q�
��0	�����2o�WG��1Pݝn�n�Չ�!������4���\3�k���YJ8h��*�������1�^�3
+��s��r�W����_K�����ı��i�+�?z+�(c��D�5 �*��(0��������7W���q׸�h�;n_���k��i�+<]&DN�ֻ�|�͏�]׾�)'��Þ�G��K��6��LPĝ�wQGD�x�k6�$������#
�(�Xu�T��G�?o���� �����2����_�i�<�&�����,�����RK�#r��X����ґ���S�uEɱ$��Ք����C&�>
�L^�V�J�ek�8iз����\|��N͕kݜ{EM����RKd����PN�Gt��V�����g୻>,1=]p����o�㌺��k��7s��瀛�����j�?PK   DU�X@��)  /   images/f58b3b66-0d3a-49e0-a328-e802f4e45778.png�{eWM�5��I�� ��w�;�a��]�kpww'@���;�>0�溟?�~��յ�ԪSGj���Qj_�q�(�p�|�@@@"  �`��롭���w�t��熀����1��
W�,��sރ�ch�!��թb���A&��A怳�>���P1��c4�{?�ԗ̈́�p�i�7�o���q��'Tj��7��+ ��x�t��5��@�4ic����}���R�&�%��_�&D�]���]f3�d�Z��4�����H�Dc��K�j���]tЋ���2������o'*�k7}���������vF��*���g�u�ҴR��FR�(��y�J.���{���>u-y)��ȕ̚���7���/��L�B^��Yz�v���~rm�$�=ھx���%����$�p�(�ێ)�b�d����RW��#|t�#ge������&$5O�v}͎��l�<��էa```v:_��(�m�Xd��!�wgKG�}p�9��q��Z����*��Qp�!S��r0���t{�M�����/*��s�OV���1����3�eȃ0 C1�H�1��Z/[,V��c���~h�~��y�o���}��!V0oڦ���\�#�<��n�����E�v4̥]���<@ �!T���x�ف&dlJà�m������b���-�Ɨ��u�(#x��)���Ŗ��7|x�Z�j�S��(u�2hU����Y��W������ݦ���Ԁ@��Ga߾�X�Qm^�{0xy���pg����w�ל���/[��cu<َi+�u"��ʨ���۳��I�#�Uc�&�[������׉������ܱr����X�rAĈw!��/��6I�˻/Ty�O�R�0�,�8*ɽM*�}�վ���?�kV4ʷ�%�Û��1��[��/uzM�g�P��_a�'y�|�1���!�cQ/ے��恑�x���w��0y���#j^�gX��n�DT}ҨL�@�"9�=H�y_`�~/*�W%�L�kH�3DB�5,�W�@?{���<��������ѻ��껀��	��/b[;��W.�܍d~UI�o�/����R��6�P�wWа,����T�^Nw�A�֪�����%����t��'7��Iy�-�r�|��cC>�܁�������k�8TZh%嘙�k�,lV3�U��{��T��}@���旜�4ӏo��g�.��Bv���sfK=s��:����ʷ���L�1����]�j���1� ��6��uj�[~|�eĔE ���^���/�O~�бd��v�z�7s�2��L��xm�$dr~�t��������L��E4O���q�~�k�9�C$�@«��
0*�9�A-p����"���A�ݻ�ޜ��۟�6�[t�s~U��q��x���}Xń��y��m2ß���É���R����[�gb$Q3�AȆb���$l��TDl��4�m���NIͰ$��te��S	�)��>�9�'���B�Ѐ��k���vgCFt-*�P�ط?eg�Y�ny���N~�
�57{zz=���a�	�ãNݧq:.�"G���-D���e��'7u�\aww���jk㷎wuj,8˚3�"�/?*K��:�%�����v�v2�1�bf(1?���4.�I"ɍǬ��^��k�N���ɢ������"�ථ�T01�Ѝ=�ꊟ��:&2��f~��P�O�Lq�?���N���r��`l�e��ܫI8�������)�,����_��K����>J��r�9Ih~yC���)!���5�н}������[����T�'�-�>*0��ʏwLx�� ���8?�|��PK��O)�I/W.�v�x;�0p�R�l˘�)ո|��,���/��'��:,�d��T������u�b��
��%Br���w?���iI��Q_bu���qՑ\�#���#��(a�t��qeg�� z��"H����l�D���b���.�ө�n��\{[A����a	{Iq&��K�vGm��c��q�h9���
j�h]��<)Iw��q�U����դ�倛j��^ ���������\���D���->�ao��'e�讛���K#��L�FPJ�p���/�_"K0v��5���h�	�80�kw��t�y�V�����U���O�Gl��t4�ʱp�ll?%�!7,5:���n�(�6�,:��F�~��%��OVfJ�z����I��P!�����'�A��F�3���촗��p�(�?T�E݅аA�F��snA�
�ϥ�=�̴�#�b�gV�-�g8����;��'*.U{q��  4E�~���N�I'���P�x��A`�*p���C���Kښ�'��O��A�/6���ކ�5�-'_dD�ۦF����Ά�()��]�KLjQ�E�~NMq* @��5���C][���pQO^x�/�-�&y	��� ���e�lYfʷ�iߝ~�k����}�6z�{t����͞ �N�qC��:;1���ަ0��)�U���vi��C�s���W�C��e�C�t�4��zp�X�_��W�����|�C���Y�å��h,q�W>x����q�������Q���Q%|u� �� �!lg]���i:���x��0�2�p��Trchuy����^@�xiy�+�Aa�N��7���]@4F�&�e��Wl��ȶvu��4��J<�_�a�n���^����h�3� V�ɏ�0����f�N���;��iu�K;~���j�۱�
���	�p�9�����Ew�'11���>{�� ����Xi��n�^^���H��3�@� `���п�jYY(��A�tޠ�������S/�:c��a�l�z9�51��ǡ	���.�ɘ23��K��~�h����~<۹��c`��.-0�`�2B��Ť��M MH�c��2�동k=��y��4ع޻Q�S &&�0����f�~�Dp79y���b�2��L<~�/״���Wz\y�-VSYؓ p��y�5�m��(�uq���{��1��c�ɓ��Oԝ��CK� �4�q�j���Jt�ru��e��c�^�Ӗ��󅤋)�����iP�rp��������Ѱ��K��9��L�����l�J��,����@j�z؀�8��)�����:����P�@��Y��+�;���?��1�p�F_�ϟX����s������>s!;�K�.��?&F2[�i&%�,ߧ��AE�o��U���n'8���?.pr|��~��"�9������Be��t�0��Is��^-�����V�k��]�������~�2����ԗ�\���I�p��Ʋ���0�_g���)�t����N��SR��O�A�O���� �A�酵B)o�&	\��ᖨ�q���?CK)f �����}�Tz�������-wfm�J�ʯ��&T{Y3�E�\r����8[�O�����:L\�A��.�
2���N�;&�i�Ut�����s�e���K��C�
B	W����n���~��NM%�����Δ	[��]DG(9��(Hs0|��T��a>����{L�d���H�ю+�S���ʅ�'$X���P��k�ζ�iS6�huI9g�TݓKև�=�w��$�o����''� �;̽��������q������أ��}�GnȨ�D���Eϭ�z$�mv��C�C�e��a.���}�î�d�"��_:|�y�,4gZ�L�1ɺ�z7P,�eT�_��h�Y��;u=�A4u�U��A����8agF��!�@�� ~7[��k!߷Qg����÷�Da?)�%�UZ���=2X��=o�5�r�+�j3y����s�$Ʈ�}��������*9��2�p�[i����~m�(���n�g��Y��v����h�T�ɔibu�3�T=}�"�MZ�:-6m�_�>G����Ↄ1�C�����Wwt�I���i��f	F��P��8��7��!z�Q��Y䖫*K�_)��z�C�r�;j��v�-�%�%�XNi=�a�[����x��Dww�Ϛ�h����Jj���hQZ�;�|����ܭY��f�
=y�ne����ֽ���X&t������.���t�@ � ,�˂�s�}M8Y���!�� �2"��>���
]��b��@�16����iE���fO��Zz��61�Dg\F��,�N@� ��)舞J�����Mm�O}ɟ�C�`�}�!�7���5it �dC�lL�$�I�@0*`Z9��2��`�x���bM�=9��m��:��?���N�X��u����Q����;�#�ï[�~#Hqi�(�O��P�w���w�����"	���W8�@P�&�u�kg���J���;�z3����{'�&.�����zT^����l2�>M����!UG7>�o_�{��r�&w��/6Ey��~��<kB���׻�N�I�p���f
�&u������C�Ǧ�;����U�1�������iDJ$�w���v!sT;K�=Տ{r���Gj�{hN����q$���ͯ��X#)aG��Gy�^��	�4 �C�	�^�X�&1�O�֫����D)�Fg����S�L!G}���ϼ(nq9�2�tR�+��eF���#؉ey>�NR��g��?��tBy�L�}�Or�:\K��t&�,GY?M[q+1�R'S�Μ�4�G�oֶ`���3����|���d�H!E�BΛ	��.������W�ɪ���!}{q?ڃ{�fl�|�J΁���e�8�ސ��ìs}J_n��R��.���ι�7r/쮎}o���=���0��B4	�
κ��ez�Pބ�O+��MMf�һ����I��3��O6����L�?fn&�ٹ�I&�)�z����= �w;zm�)�'��'|�����\���~ݚ��������>�� �=����L�o��ę�r��{�#½�o�wm�?^���]�s-7��0�B�����$���\�D�O�c������&yG˓���43�6Fcq��dUK�:4����Z�X���(��A����wā���#H2��BLΔ� �u~� .N9w������o�^�u2i�x�5�5��w��<ay4�˳HI�/��y��X�׏�II�D,���Hė�>����S�����S�_䬺i_��'a�e׎3��f�֫G	�?Kо0l$�2�4��,���wItN��f��s]w�=ےqh����o��x�@�|Q2CX0��*o(��r_^Q��ֶ����2vf�=�6hu�B�M���U��;=���s���~	��z8�B��sJ��W��w�Db%�������{��2m�ݗK��w���R����&Q,����U�UL^|�Z�$�%���d�GҫwIC���.����~u=2jc-�e-�U"�mo���9����}?�Y5��8�K��~��b��(dk���#&؉�A2+��4�2��&�(p#�u���^b��}Vt=9�M�q;�u�����S4�9X���N�A�ӗ��(x,'�.��r�j���n�\��K�MI�T�W��2�����u��uP�l�����ّl	K���a҄X� Oc%%�Ж3���J�Sd����R��Yp0�0�tXF����0E�Z�T����� ���#-�B-F�܆�?�]�<�K����o�	�$-3</M�_�N�f̊��~�x��)�Q�En��k���?ĥ9�ZY����x����Ìi�{��d�W2O&E��_���'*�N�
6�+<�.R���S�^�G͊o&BT�7���3K�����ݍ�o�0~�0���Vd���48B�Df8����ƾ��Ѻ�ʑ|r~'�"Bm����wK�lN��b�-�37��:�������h:`h�t�2}���;��-�)
6}h5���LY�� ̓^Mj{����6}�:韬�sX��е���'�W�P�g
�l��LI��g"�P<A�9�a#�w�S|��1�H�8@_�����fP��qQB<��6��
��T��I�as��!S�����S#l��}�t������P�a�蔏���un�(-@��{XV�J�@="��u9�f��6]�8c�π�n�1mڒ����d]�^�h��c�M�֤�8�f y��} ��Q	���x�^�;۸���L��ܢ��:f�$/�駭��B��,��/!��g�cۓ7���:	�%~ �J�O?��������X�sG�</W��Š���f"�
�u�t�fC�s�������4�;tڇ	�c���;B�dF��3F��
s�U���o�KE}�|�	=��9�&�Hs��|�C)���	c��*�n^� �S�y6A��/$=�N�1&K��i0�h����ߩQ��L�\�%ޑ�I�u+'���U�U���/�A/3� :Z�AY#C�{��:M%�5�-�2���h`���B���fϩ,�f�K�� Dc���	W�@'B$7i���#�yDh��IoFb�&��_B�����4�� �#�\c�aA.�%��ھn޷��UjU	,C��^��=��EU�($bP��rq�℈�?���BT�Mm�)�Gj�d��z�㦨�OzG��|��U�}�т� �.����������wb���ٙC,ddD$�hQ���q#�� :�9�1=#�Ȑ�X��Ǵűo����B����v�X����S%S��!�g�VrLo9��/��:}s���~�<���j��h�`D=W�g�������|~\��<va���|?�=�ď��٬<
?�vJ���M�C�
%�� �T�h���>�7~�*�į����ȵ�H($�
�Zn���E��v��g[�?Ĥ:¥L{�Af�b%*�����3T������G�i
ߘ�jih���&��xY�O��fB�,	n*�×}��?��V��NeV̛ X�)�S�';*:�2<8B���:&5��їf+�N����=�V���2��/�)~Չo�u�&��N���v�y*�'����&����޽�\}��O��3�ןf]@��o�VA@�<P��]�:P��1W=���k
9�����5�o���~���b��J������qpW^�W����q3D��GX�a
���9����������d�o�S-|�>KU�@/�J�t���������x��
����shu��}�h���_�����|fv��o�M���I�>SD�K��/]�P|w��=�	7U�2��mv���٢�I�D~���z}��	����g̻�a�&zF�#u�F:��Ʀ�<CHJ�����m�{�|Э��Y�f10z��W+��C�]�Qz@R'a��]/	Q�O�����Gv�k�L~�x�Jn��ʻ�[��y���bI��H�lۗ�8)ώFnE�P�U�[cW��q�y�t��S��9�"�
|X��:[��J�������O�4���d�m�7�q\K�,"y�=�T��	C��'��c�J��ʕ$�&���į��#����1#X����p�E�.Mw].�K����1���	@���87�N�'Lw!6�ۀ�5���=�?D	��F�~�	ن�y���<9f[T�	1+�b+8�m�R�JO��Ũµ��Bgw��?�F*�.\��$�x_#���7��;Yn3�j'�����=]&϶��D��ID�x��>k�7�_c |af*PF!@7S�� @��o��]}i��f?�"x4�IwA7�{y���nwȆ�4�> �.Io�&�p���kަӢ�֌2VبXݘM����X qJ������Z��=1���q/g*0{YY����;��d<�/�����_R���*�[��Vݤ�*�ڜ�fS��O�ʲ1�)N�CɎ�'�������5�bc�s��ID�Ή	�N�u�\����7S�kM�"&\��2ԥ�^:�s��b�#�po"�V'-#������Xkz��^>������FR��Ν&��v� Ix7���^�Cf�� �H����|{�	�Ce2&�?��׵��l9�^"~��o7���C���/K��~O�w�&G/��qvm��(�&uv����7{��Y|3n<�#�Ɂ�Kl������v�X���(��{��!0�2qƪ��\�C��D	f�n��_4����Gx���^&���|"�V�-�N�����/1v}ŕ�����oӉk�]Z�4����_��t�}J&��MP�G�h�	�+��4O����Zy��m����[�^�RXi7kz9��\$v��V-�>�_������Λhp(��:;�{9q]sl��wy���x�	q}���EGA��+Sͫ͒D����A�Y��oG��G5T��E�]-��D�ep/CX�H�QY6��0�ة��hK$���J��N�Ã�C��k7���ON@���,2����l�r�����p-�'J�\���9�����a��e.
B5I���â�s����.*����=�K�?��4�f;�:�׀��B��B�aJ����1V�O�)��/�E��Fmcڟ��}��_��t�l�2��.����1��g������6R�������lN2,8�
�]�S�����S�}U�@X��Ɔ�Mve;��a�0
$��P)}��7#.�T��G\��lp]	>����%t.����V���΍%+[J� �D��h�li��z�X�� nw?�x@%�>JY�x��h�VP��l�Sw~Eji��u����|�M�6���j�^�n�JH�ؿ��dbMߋ�̬�����F��U�!�k\��O	˴�͌7T����r&�m10ͬ�:�j�����ז3fU��Ѳ��W����������E HRBt�U�(�}f!�JBN�,km΂L���HVӦxG 8t���h:�A� /ɒODO;���;�zo�;".�G�,W����%�D:�C1C�5Ŀ@������z)�Ɍ�#�2���OR*dҞ:����ıd�b����t�q���c�׏��q�s�{��RQ��+�ж�mi��s	�l!���UͿ�!�
���)�;�;��Y
c�)�PCp��N�G�_�E;Wh�̲e��	���̲f���56�eV%���e1�~숆�գ��[�+�������R��h��R'��F&��	�@��8�P�'H��E��KX��G"rr�[ZHK�G)�c6R2���=n:�HU�@6��{Q�f�aAb���<��װY�O�}Q6�w*���3��#�����I?I�f��>�%&>4��y� ���VrCｰZe�|x���'Wj��i�o8��e���V��2h}���=�)O�Qe�F2�!�45�L�4ՖuVj�a쫓ρ��j�+$���L�����BU�{�^���T�� :��vYI���
-str�gv�B{t,����kk3�hƃ/�I�'�_%߿��j�v�M 3�ѓOM��D�%�͸N�������z�MD��+���z�@�wL�5t2��_~�c�E�7��G>�w'*3\5�kImt��m���~Oq(^�˘��W¤�z��%7���C;�j����p���v��^N7	a�cz��u�o�j���'a�$��%�7����fQE	6c�c��|Π��|��&� LD\������Pu53asE���z�[_�&�W�@i��D�%���Q��kA�_�4m\��T E��3:���ÄGZ	�@E�YdF���-��>?s�Iz��b��m8�#C[�-�{�뢢!t��!���R����g�1�z��E\���Qly��1sF�;/
l2��g�(e����2`�����H�Bl/!� ��ޏ��ǘ����M�c,W�|��8d0+vP�]$B�v"��GO�����+E�a&$���ћ�P:�>K�P2kŖj��0ߘi������L��o��4�Y{y^t�<6:�V��\�{�}9I~@`��;5�W���o���j�9�ѩ�Q��t���]���k��ΐ�M�7�D�_8�<�C%�[<2��� q�J��ڂ'�B&܅1{�h�����pg�-�^�Z�����*bA�ʭ
#>���+��Bn��d�bksx��x�#}\֜q����|m~�:��'U���A�V-���8=�P*���]	��Є{��9p��Ɵ\�m�ی����o����|{x�[�h����k:�h�f6�>߂����j����<�'�(k�p4��V�I+�$���L��K�5ʿ	��J��l4���t:e��<�9�PU6D\�j��m?[nNp��)�7��.��쑙Q ��uA0��H�Lm��P�ݰ`�1�ixʧS���\a�Y� �~����i����.������|�ɜ��V� �tJvLv=rq�EZ�0+�R�b�nE�G��S+o�V��)-��жx'W~�>3�_[�x�����}�}�z~�ʃ�cQ�C¤��-	 �"$��"��5h���K����g�k�e�$Cjk*�XE}�>�~����וVBVk��'UR>�S����r6����8u3�p���FM}�ԟd���d�n�m?vR�ܼ;�?�~!�l�9�������Ti$�	�vp�}�����>�CөP`�^��,��]�&=5h~�O�{G�O����[�$�G�r������:7Rv�����IF^���9%�L�;���l���&�z�0,�Y��-S:�$���f�	9�)X����8_������O����9�O�k�塩\S�m���B�+X�9�ylI0k�����C�1{�^�� ���-4�8[��8�5N���I^J6sA����ʦ����j�QY������硖�k���M�(���_/uu$#]@�>�$�!�!����Ea��=����fw�>H3�94�Q�]!g3v6*݊4������ǥ)����t��T�_�P���6��~�a.���7",�U�K:�|/���βڶ��]�y�}*�?P��*�~_1�y�.�<���%�L=�-���X���>Ҷ��*M=9��P��od����ck%��x}�ȒMP�I�]	��1mS5�Ҧڝ5O�`L�@卬F�
�%�����7+Pۣk��I��,�G{4BI�0�1�֍�.�K��~��h0�4�E���;˺�~�{����,S�Ѵ��i��=���.%��o�˹�A 6��Z펩��Í�ݿ[�q���9�$M��<q侺ň�����+���������=ʐz~Ffu�X�|�?��}o��K�!p0���ur���8�lD��g�T�>�P7�����a�"3d�3{�
g�������J��%�����|�_#��N������f�j�TO��9=+qT�6�#�L��vf?Rk��|��g���qm������O{�֦<���K�ڝ�E������(u��տd�!�ӗ�A�vi�d݇����f���i7��тG��C���eCX0�h݀��A����'^X����'\�eP+�θz��J��A7�K� u����S~�Z4)��p�W6 �����$�+p�c����`&X��8Q�p��w����Ϸ䠊9�6���A�H�ӗ�u�pV���*}���F���x'�ssd�����1c���{�L�z��R"��o?E}pA����򩓲��Cʜ7���*G_���cv��U%[:٣����|��&��y�|����C�w��fv~]��__�F7H0���$��p<^$��E[BM8�NEG^&�ht.�C$�Q���l�uo�޺��`�4iM�w�q�j���cN9w�5u<ǹd'Y:��n�����.�m~�}S�֥���������x5S�-K��y�����5]G�_�R�-��x`P�8�v�(O�>�n�ݣ,T�XQ����w��������� yR"Y�#l5��`_��ݍغ�G!��f߅�jV��+�����ƴЅ�����
����=��޸ �*
Rj:m�z��>�XS���=:��uy��}F (@�ɽ �X}���p�&Ϩ-��a~'��J�'�:�\}NP�U�&ֽ�m6�n9B�����Z��+�V�[�=���:&���H����ʄ����wR--VX'����kT�g/S��*9 ��T�x�r�L�����J����#v�j15l��H��`����07��gQ-!���@}U��#ƽdL�6Ά��
Ȇ5��?�k�2C�r\`q՗]��b�w���t���yb�h�&`�!�+��k0x�í�ϛ���J�{[K�x�(u�J�Q���j�8q��j��@]"���z�8e�i!�#�Y�Y�1[C�u(��| WuFR��}�S�-�ƹ�0���Q���.�6wm[w$��Z��C7FMЙ���o���ZTnSfv�-a��i\7�φ��_�v��i�u,�eV�;�'ᶔ��B�	��s�a��5g����'|����%���2��\1v�Xk��_G��!��a��H�`����*�41`�~�u���cɈ��t<�	�b����a���0�$��e'1ί���e��c���
���fjg�*�c-z���m���ٚ�����a�fV��ߏ埞�7��-�cfN ���ˊ
��C�+��a��Ѧ��#���a:=i���ݦ]�W�ú�{K6����*�%��d���.�7�y3����-�ʸ����G*��N�Ѳ^�����}L�[��
H�9e���"#Z<��
�F9�6�T�B�ix��P�_�3�̪���W�f1[(��O�|�S����|=�$���b��X��٠�f���:{��J�p��j~��,��-ST�z
=C���+��}�?����X��-�H�k�~�}��XD:I��
�q�h��Dj9�+#D��Z83��På��{��K�?@݂�uq���Tȟ<���J9�!l��|�3#́T�T N_����"�4?���i������0���`����1�n�=�����r�(j�!H^�wp�e�<���\����haBxPXFiY%�Sgd�����f�*�ZH��ɩ2����tƩ�*�(RU+q�h��z��h��/�)ݳ�P�c�SPs�H6���i31�~42�x�Of��l\,���\���x}Y��>9=q�ґS��U�.����<jK�l���l1�#�������m̲�����X��u��Ē�)'�Y��G��}�e�����ū�b�3���n��o�\�G�wį�/m^��P0n�ө\��r�(/~�=4,��.�姚�LCn7AHB�٫~�#�y��cl�qt�*����ApCZS��.fe�s�6������{��BO�<ae:6텖S��:��N��.�Z:0�ͣ������o�(O�����'��f�y"��8���M��q�U�<X�^���>�!R��q��<������z�V�2"���s0�_�5E�HJ��ʿ���P�,5O�!��1��X��7Fq��̔$��j3��w� ���k��[
7��<�E�Ӣ��~��x�B
j�y�I�.yIl��}�-ɌNR�?�$�
�����&LC�DfP��R��J���݆�׈O���Ά��/���,[k�R�yEaQ����3[Ҕ�ڪ�B�l%n�k���@�K��fT�
��ٗ5G,H�ߴ�6r4�id�LB�O�[�j.��e>��f{ġ���@�Ñ$����'���䱳�yl�sZY5��s���5����k���7{� �c�Dqn�C'�q���Љ��S+)1�I&�4W����+u�8D���w�ʴ�s4�Dse���;tQω�{!H��$�����n��P\��n�y�m?���Z.�
5���%���+������/�"Q����K�K';�0+�O_���fpm�ֶ蚾C[%X�Fǳ�	��k��p��/ 5���Ge�K�;\�R�+��2)Ʌb�S��&�kS��R��%>Y�'�M������"��gֲ�����j,���<�K�p���Lz?���(�h���p��X���[zeON��B���J���qSZ%�;/SSr�A��RO�>�g%*V�9K!�����,�M���F�� �ね���ѱ০8��r��wa��'g'���km����G\�Z�Y3:��#�Mp��I��)V�f�֨���ˏ6�z�<#Y+�3�=Z U��Wں��-2⺃��>Ur��|֩^n��n'�Io��D%	Nvr���f2᪣�L�!JÞ���7����[����̖�����SL��tGy��i~�Et��TB6��O�Bz�-V*�A��o�Nb#W��J�,�W;�EZ�h�~-��:��
�H9��i|�
��󝾶Lw(a�x��ZG�(.��<� _�;dּ�5<�?C6���[�D~p��ep"P���4\a<�|�E4��CLT�Gz���P����6~)5�^R��4+�{Oc�m!��U@��s��~#���Ygw�Q:{ԄDA�Hǔj��`�l���m�z�T���^������(��y��yo9(^<iJؠ�X�D�H��~3{�Ze�hz�A/��ܬ&�L� �q�} �#j���U�ea����m�~c��J���l�
�R��3U{��a@ej������7��U����~kz�j���vi��&�h胃F��%=��o�ETYB��&F��l.<?�-I3�t�'aV�D�^�$�~ř����闧U�p�$�d}!q>ah�Ă��~t0�jn����#��)��Uqs���B�����	RH�	Z [��������U�;Lq�t#�*��9�#gCp�mX�B��bj�U4��ݏgY��,�}PZ+���OZ�YMh�l�dH���c1�]�tP-����
�jQ JAq8��|��Ҡzc�Gh#��p|����2�b���QI��H���;
W����	[�e���ALK-є��|�L8Aqrp��s岎z�B��5�Q��0�b·��5�X�H��w�~f� �i�p�Y�~�.ஊEH�4�/}�J�hu�[��1��k/o��|�ߊ�d�cf�AcpWq�M��oJJH���t~u(]�ݚ��F:VV����GL����4��f��'�������G(=Wa��?��)7���`{��P��s5b@ɠ�4	�03��+�߁�pߔWH��^�M%A$^9�>�L�o�NEt8A+�=�?1M�}a���V����ϥ���l�'@a�dI#����h!�H?�M�i��Y��Q�m�y��Sx�%պߙ�!�G��0m���ɓ(�B�n:#	ڹG��$γ q+�x�Ɋ[dO
�)�@y�>yS�-8.:�=�W4�k>�f&NWtO`�^�57H6f25E���vi��4���W��Th��� ���eۣ�ub��h��U�7V�7j��kc�{u��M^Ou����p��}�S�t��KSf�`+�5K�F0��G�-��ݴ%q����2�P��I�D�����-��?�i�j��"�lqln/aQr��[���]�d�XL�B�O�H�F��ڽ�ϣI~�<�H�8�q�9w����-pcRފo�5W�����6����y�_������yhiu/�pS�(WQ!�O��hn�@���r�|�U�Vfٛ��!�㵪�R�+_���6E�f"8�i�)bR�w�p��X�rҹ4�؋�t�vDU}����ΆCo��#���X:#9�.�%��7!��W�d�q�Y�5v[&!�/6�a���&�}Me���5��\�a�$�K3�=�Z��K�y|	�x)v��3h
I�k�8[���CY�9�"-��b��ʲ�8�!�[�ed�Ρ?[��m�gAX��Q_2!�2]+�*�^���_61��ΐ����F���c]׽�J0��;ad��n��|43X�����?g�/r��h�?I�tf���X�f��N7�i���:4�շ���T9�Tɝ�l	�%��5�J�@ա2Yg�t�<ԕL��KO��W��|І"Q��[97�b�;V��K��F�]���}9~��-�
E�AЅ8���e`���5�K�5T�-�J
�� ]��wE���d'�X��Y�{L�Ͻ�/��pd��Х7��ofM�$��n7�n��ƒ�P���z���6kjMx�>!�O��G����D�����do�� �����}v�zﺩᩋ	���=�05s�T8��x���T%`������f�P�F���1���i%�˥�9�`\�&�����Y�s����S�l���k�t�����|rZ����$7���"���C ��	�]ωs+5Nf����0�?t�k:�V�@j5��泥������hƄ��m�"ywc������N+�wa�,��6�9c�%��J�Q ��qx�e	�;x5��������HB�	���$��#*����v�յ�?9"M(��DV~��Z������N�^|�k�S�B���Ch�0�'�	����ŕn�dc|��`@����=���p�NkWm���F+ox�l���@����U=�}�Q�7�I<�`2��� ΑI�R�e���L�J���gA�^��-�ˆ4n��O)@Y.���߹�*���?nnl.���,?w{�e9xn�c�#�g2!�����ԇ�p����� ���֊g�n6jg�ݤ�D��w�k����<B�n�w��ۣb�=��K����O^X���+�.�L͗SOYf�j) �"(�����3��_����L>t��aݭ@����_��X��?�Vv��Y� �\r�B=��u��7+_a�\6�Z����oy�{߫��I�r�����{�<��	A^h�ha��,9Nλ�U��̳����m��fx�^].�`kq�{��y�{6��	���4�!��`��nيSe剧� ����|ꩧ�� ��yh����Zy��U�c2���7�?�,Y�D�z��������؈�E���}W�k��rQ�Ni�\���0����faiٿ�[3xӞm<W����v�1Md�̦$b��6Ԧ @������ܢ{d��sn��`�{3���fdS���s�|<�	�,���eB���mA�&)�x.6*aͨh�����Z���7�n	c
@םq��N*��e��?��I������#��r���m��B%��B���=�a^LJ�l �!����ݽ]
���B\�L�=���fM��j�a�[&˫/�B^{����PA��)�����G��C�ۨO��c��>�6���+L�I'��e���Ym���������a޹���y�0  pL&�(�ʠ0���c��]��ʕ��l�/Z�$�d���+�/��dD.�u{�r��%=��q�O��g�cNF���C悈�2��m���0.S�k�<��s+M�j���)`�`�N2V�"�9Y�Ƶ&Ș]0�7������6�8�E�(x�
�;��m��� �� �XS������/lIg��m���e}gW�(J-f�H�`�H�b��@�iZZ͝�/�5����>�Y�H�U�fLozӛ�G?����|\(8�:H��A�� 
a�1΁�q����{�9���uP�9|ͱ�&n3�!���VѶp,�t��Y|��CK�a����I���h#�YP+�y�+����ʍ���ovъ7�&Յp�={�Q�^�8�S
}�R�`q[�V[�y� �nb�?@��o���<�DW�[锉u��D+�� �mj�Ԩ)Ad�\ 2K�K!�j�Ԩ�ٓ�������S��B���jx>�R�pKoP����s][n����砐!S���r��D%��Z&ǘc;�)hf'�E%�S�;+0"���9���)Ӎ��Sk9�N)�ӎ[_c>3 �$��U�Vi�}��>4z0v|��|@���AK��xZ�ZV¬'Xp��M$��Z����Wf�c�!4�
���`�3�`��orB���I� C kD��=��D�Z]0�0AH�:��4%E��9��&S���q�>���Ae��4Z�ʲ����{��[�Fv��l62�X�ڪڭ��S��؅3�5�	�^1�`Xd�7k��[���1���9q���q�ݾ
��ϸ �}n�}U�c���?X}�|l`ι+�"�u�jSxP萑��\�����cxM*9n\�֔ƋB�D���*�V�}�>G���(u��.>$UyAY3߳f��x�L��@�(iM�V�y��k���Jv��M��.�}�z�ɚ�w/��:a�����^˶`�c}2>B%�c��H�A�������<hR�YK���Cca�F���# Ԣ�_e ��&:M^jVdH�	]F�����'�9�	�&7L=������L�Z�ٔ�4�8���2y��j,�}{wjuC<������c�\Ư��76��zfI�C�ɝ��(�x97�;6���q��Ժ����2p������$L�q��]?�мO��.�A���i�3��j�T�sq� 7��bl���3�q�C����z�TɨR0x��n@V�&ok����3g��!FѪX�3\: d�gRz���ף��F�fQ	����Ý��|Í�p쨔a����G`n�t���o� �7T.�4ak���ΑF��e5@�'��H0X,$�KޠT.EL<ה�����ӛYtA�ܰ*� � ��P�Z�|h2�Ajl�ri�R��Ak��1Q�@��}�?]#��
�4�kt��*8��s5�cw�i����� ������OF�Vo�68:��}��Q%V��;wFnBׂ��B�G�w�n �V�{b����.��2=� \�َ߃\��gD	�p=h�(3 !F��Z0xKbk� �lT�G�؏�DH2/�����*3�Y�ZdAֱ�����ڗ��S�k�PR%ݳRƒ���c�*@��芳�����z�5:�pc�0���G,�`����	�*�q�tsj6oh�R����M�h��z47DD��0Ml�FZ�į� D���8��R��@.�!���q=�H͎.�Lʞ��&C��v,۰)ߨ\�ճ�`��i��/2�t�X&<����oW�4炕S]�>��=�c7�t�n>7�]����;2N0�~UPD���
��Z�h�1F�}�_q����~��������8'��abS��x�-��d<\fH0��,@�0���	����������߯y�k���>C�_���� � 0@�l��Z/A��6��BU�޾^�_ 6
����V��,4�?~��(yYM��֏����
E9w��7ܠ�?ʺCQ���
~���댖�Zfx��s�X��`L`���q�����f��v����L��f
_A��R��B��G퐈�������Zh��k�>{����]��ɧVK�*}���Z�@�YlQ�ޫ�G�;�O"+-��.4-)��) Z�T@W��v�8�Mr�>��`=@��&eB	���q�\��K�.�x7(��+�g���!M����`�{隵�ۼy�BfP���KK��up,�{�'��\ (`�x�5e�b��!��KZT�:��"����F��{����u��S�į�_��g�2�W���rkn�"�g̷E���ݣgq������ *JVٲ�����B�yC)g�E8�T�xp��+�d�a׭��v��B��1*M �����#�礹Z�;q 2w�(�M��Z��+�B�ߥ~!��ν��COjUO�=��%��G�n]���f�$5Ϗ�:�7k�'�#�%������_Z�{��H����6͋[eQk����܋-��$޿�����w߭��:9������&����`ʌS0���Ƞ/��zX8�t� ��f�ƅ@n^������,�×���~���Gq,�����gsv��p<~ñ� �|�I٢�O3v��B��(@�U�u��SOJ�-Z�y��ǩ+4O�e�&��0 o�O����[��`�"7�H�����q�� ���`��S
�M�Av5|��r%u܅� #�@�Ƥ�ZRm��=��<���mL�Nm6�|����n��֐�^2�-���������� ���F�]�IYa��H.0B��B7m,%-�e6=��BW@b79j-6�4��z}�[%�;4�@�k~������� � ���C�	\�0?���� ���r���eP��Q?� 7�k�cG��!�tAo��袱L�U��k|�\U$��2o�+�j�{�N�/�F���	_���%t�Kk	h�����0��ZP�h�q�k�`b"������Bak��?��gRҹq!3�B���es��@n"�L��Ԉ�v�b��ohz����ק@�����\��B���6��w�N��]Q]=V`�B�n����_ށcC��9� ���h���
 �#H���g~�_����0��`&8�����Dt��."ąC2�ߏ�i�L}7�׍Q�� ��pqshE0Ǆ�D�ؖ��h}�0O�/QP�s��5�ǔn�1�u(��^`��5Np�:N��3Q �|}�b�� ǂ�(c@&<��ts<��606��/Aᅟ���TF9wno�C�	����΀�3qӻAN,.|�=>mdsp��:l���.�:V����W얖f�,GG��� �y
}eim�&۷�UV�Ug��:�4�7�X&b�� �(�_{0&OA@���,��l���Q�%��5]j�86;|��3�b��,>�8�b�q-�tuv�0b�<|��l:Zp���5>��I���q< ��d�8����?�=��83�)p4���\�ŭT�ZXcO������9{Y�v=���B9�bE]�%-����C�K_��&��Q����z�9@�C_|����q��P�y�_��7���+����omrq� 6}�4��F.$���k��(���M��f����Ѓ!U�[�R�5&j�4�=X2]ʅ�m�e���Z�X��*�Mii$��w!c���3�ʶ�.���w�[�����I.y�7F�}��`�6���\p��Ua�a��
��[�S&������`� O?1�y�d�T�������k}�k�q�x@�L���7D���Xo�jH� ��J�lI��1
$�V��gl �#Z�`�e,�*af}oݺMv��"�]����݃]M�R���e
J�) "���泮C?���T{���\��J�Pֿ���u��O�r����:��?����#C���T~�\<.' ���+������E�z(��ڵO�=��J��\�Y�[���
T�D�K��֠�. ]L��,uiycMsHd��w�� ���|�)2�?h���oFv	�
����;������#D�v�✘&�����*�87�F���:��lὕ����c�7�	��V!MW_}�Z@���q#c���z�*���O�T�&ċ�̃���@ny�������2�I������c��@c?[��{�V�\�x�\|�%�kj�b����Ui��|�H�P�����B?U�NGx���=��c*�+7��E�h���Z�J���*���\S-����~�'���#��-�j���6Lm�I\<�\��bc�*	Q��N^5��Æ-Is>-My�8У�/� �V�`���m���O���>�}AK��A�:܅ձ����/��PD;L���,Y�9���
,;�5`l4�/���'�|R��c�6���~����y�E�
w\��eR�V���$��K$O�m�����b��\Q��н�w�Cq�����d\L�" =�� �YXXn�9 ��3�0��k����.����|�[���Q������/̾��%G��_)�TE B�GU�T�E:���}�,Eb�=,��P{8�󬲩��la78�Y��M֢�2���������9V˼c�����C<(�^\�%f��N�+t(�2���ɠ���'/��n��C#hmn��^q��^li�k�n)4o�0P<�}�4����Ȏ۴�+�}%�fWC<��(��ۆ�]�2e_q^%b$�p���!�l�fq��$����+��@Ҿ�V�,i�(�b�����j�Ę��4��e�Wv#J�>�'Y� D_4QR`~``�`R[��8n�����׍��w6�p0OM�:��A��q5z� 6e.�U�,m����_�B	��Gg6�j6o�$�=�Z�Ο#���&2}�4Y�dQ�L?%��T��L�h j瀝~�{ߋ~�~�!��@/������#Z�T\p�w����)p\���I^6cW������^�sF;���(H���=��@Qjn�*�Y.��1�A����\�W��@AT ��c2�xr�)��+�kk�Ұ.1��vݻX3hԂns���u���e,�>���eR��C�\�Z]WPf�e3[m�\J�+��P�y�3���>ʲk�G��k��FN;����rQ��:tĚ>}�E\��`B_w�uZ��6�x �IiYpBt�d�1���k}�|��u1V�}�g2ZO�%b�� #�����;8��e��k��$�*d� l2�M��%�nj�����K�:JD��&r���w,Ǎ�!��H����(p�(�+������[*J�P��x�jts@ns<#��<�PD����V	�נ["���-�� ���};d�]j�s6�f	޳��y�	ZP�J���E(8� %��#d�z��}l)��ZO�ׁ9����#����R���׀򁜌׾�r��F��۩ �fË�v���5�'g�q��6�w���$�,��Ϳ.��g��d�Ye��^q��r���F[��"۷o���{��Ӻ�ʁv�9��Ur��ʹ|����>�#��b�]�9>Wl�!�/#ӧ��Ν�d���֔kֆ�U�Zj)ؚ'E���i2�Qb�fj�����H��"p\+����S�fi����X\+�����x��P
���j��j����V���g���XC
V5o֕"���	"���ȃ+}��``��`~Gȧk}��4�9V����B��92T�tQ�X�:��/L�4n乂����VY|�rm�R�x�W�\�I���S5��dI7K���h������_��_���B����&�ʤߞ�EZiHXl��񤣳W�|�qy�чuMa.Qtn���SVi>;���<���Rr�D�b��{�?���̀	[�p��y�*-�Ma��r�}��R� K�_�Z@�`�c`����m�������vO �#,5Lm�f=�7����yg�M2w�B�>m���K��κ��ul]r��À�ϩ�9�?�I�]�>lb�3w�2a$��Dl����1��A7���k-���R��V?��ƅ��!_C��HVz�pu\���� �u�� (�6N�r7�}���h�=��w�c=:�>6n�[9�*���g�]��D�j��=e��*֌��ڦʱ�N5V�d����J;kR�γ��E���S�yGa@X���1�p��1c��-�o�p1G�c��Ռ���J�7��=&;w�0����m�7���O?a��.9�3����SČ`Yt�t`�;���h[�dB��x�J�	�	�g�9�x꼱
:�&�+�}�fО1��+{�w�r�u��	?�St1���2W�[���Ѩ��|�fvw�����d��=�չG{���,r4}�ثha�r��c��m�c�	ƅ&:�h0����5p��D0����̰9Yր��A."��&�t3��Aӊ�@�B��tx0��	 ^�&�L
�=Ρn?Ϗ����ʡ�?�!f{��E�!KL@`�
�O�����H#h��$Jh(ˉ��D3
Z���Ǟ���}.��1��P֘@���f�L6L�j�)����K�h)���z��%��,�[�����1A�Cq<}�c�X���Y��D�pЧ7(w˾����m�Q�ɓ��W6��QZ2���+=����+.����Y�Dݍ��)�!.���'jIg뭫C�M�F�L: l�s�����)��z�̝�n&�7Z��P�����}���
�Ǥ��؄��N�5�&tr��sf1���H���0�L�f�I/V ��u� ��0=TJD�K�KA������e�����S2�K�/� ����7���������N8A��N���ʏ�# ������=�I�e�9I��C����o~3��Z|X�lr������k����w�|��%�i�����uP@Q,��}-�u���J�{�U� x=�����X�F(V+���f�K-�ַ�U_�������{J
�����Z���:�%e��������M4_~oo�TM���^������[.X,��:S�S((�z���@�Ρиg�A�HPH\�S�LW�	S)϶jKy%�:��h�6�J�5��.D�{dR�$ٵ��M���Z%69zw��t�x��~�^�E����NYֲ��im�I.m��r���E�R)!���o#��Z! �XOl6�Q�o�� >C\4�0@�.�G�+��:0Y h���+TS���������|�Ҙ6�]���2�pʤ�
�۷�h�}e�+�����w�B����5�gd)
�qpO`T \�)��������5F�s�O�	0B������
��A�J����j��]pġ���d�_��v�/�˥�2o�!�cm��P4?�s`�̜�D�F�+�i�T���s���SU�?.�7˖/���g�8m�Ƿ��-:�_��Wt�1Gl��?�vwȚ'�ŋ�Ȭ��e�_�4���^�3�=�roi��Ï<(�/]a�grdMn޼�Go�3͢��2P��ф3ƎZ��93�6��l�~�L�fi�e5��VnՒE�Ф#���7��C��\D�?�zܐk-mi���'�o�M�ךg(X �{��- �?c�\'1���h7!���nA5$>Aಅ#}���c������������$8�52W\��MX�((x#@��+��2�� 0Pi��#-���&����wn� �k��q����_/pK��ѳ�>��G�"�@�k%!��6r��D:�@J"�@a�u���%+��_���eS����e��Ge�	�$�d�~�(�j�%~�C!¼3~��}׮
���AX������K��	�פ�:��;�aƻ��ת������̄�
%��n6s>$
�:�q0~�q��=p��A�ɕ�If�E��[�[��,��#BX��Q}���m��_�����;�!g��)���m�ҴԴ�=#T����O�T4,�(�,��%}蔟Ua�����C��J��)*:�p(n������}6wN�4vb��2x���، ��]�	�bW��0��i��������<t���w��C����Ѳ�𾨀pL�}���;��#�{�6D.�����8�pq���RPQ���g�\7���<����p2T#�3�M�6���}u�jv���X�3��N�9k��q����[Rf���=���c�v��U]�{h��Gy$Z[ �0���]�7�e�+����	q,V�| N��b��?�y]������Z�{���}��0���o1������f5�b��S9�M[,9
Be��S�<����� �!͙��f�h�A�*�XHnh
�|.�Bɨܶm՘�״��V|iknU���#!�h��Y��|S����3���G�K%V�g�?d.�r|>��*�4�[4�-pr5f�,1=O&��{@.�хK�̏�w�%�(-���Hp��ܠ,����0��ɀ�c�2l�QQ�x�i�1�D.ѺaN��=����C#�K����@ �4N�ux2Z�1�^��a�a_@1*h�W6g��t^�����+�j6����X`�yͫ��y��A���,�����
���w��	�
����
�2u�qъ�eZ�Q���Y�ip9�I+��9s��!<�2�u�憛��?1��PD7 &�����6���=Ř�U��U4@5%��)��}$PuHW_��Ɛ��877]�(I�m5�!x-$
�ǲ�O|���1Y��t����b�5�͒�޽)�z�t#Д�2�`���M.�����9�x�.��ޣ�&q3MyW�e��������Em��Bf��� *�-��
>gv���;&�1a�P@���ǭ��<�D����/>���?W耈v"S#�g���
5�1�C94���*a�J���߾T��7J��Հn�Q�̝ky�����29mʲn��޿�Eo�EF!	�f�z���h�Y�e]��.C�M�k>���=�ܣ�/�ti	`<�Z'ˌYs/i��gsm��t�î����Im�F �x��3T �,��6�����z��?���v����}{�q�d�tvwȹ�](k_xFt���KS�h�d]f�m�$9jANҹ=2g^��d��ps�Իꪫ���D �����N����(&p<nb��&�M�����}��K�Lj��+����V/�@$bf����"�m�X�~4�u�nj�.4�ڸ���.��L.�P]+­�J���&�1^� �fܺ��5;W��o���� �����(���$өU7&�rqc�u9NC) |>�y\F��	��0Ǆ��Ұc^��B���R���9�|Æ��q`�с���d��^[�Y��ß� �$�L�9��0!�hˈ��4)�w�F�v�ؿ���kUY�AY�9>�' �~��� . ���K˖� [�m��[v(P��y��PpSk��O�5O����j��=,��>'�]���R��~0A�>���<����<��cr��UƼ�&}=�̝�H6o�&���/�*2�\�Yc�Z�ȢE��Y�\����{�N,��/~13�.��ԟl
bLH���vh@��~.:5+添d�ֵB�O�u�����tQ�j!�]MS���tv�� ���ʨ�[��M�'s��7�C�k���A.f�ǻ�DfF�h�E�Z_�8�v���d�|>���j����
@WP��Mܪ�'�I���q��߱E�`;�]��q�R�G�%�g�[!�E*���3{��s�z��^:s)�?��ޒ���<u�t	�e��
��ɀ��Lׅ�Ak,��)Dρ����>��ʧ>�)��~����H�s݊ p}�֚�|�lE�tv�ɶ[e���77	�VI{n4�Q���'���3t��ث(���r��R��_S�!.@�M�[o�뮽Fʥ@��Y �k!V�?��J\$U͘1K��XN9m�6�����[�zu���O�G`����Gsh	`��>�� ��!& �VS{��r�@�y���ӹ_U�\�G�v�����d�
4��2|�h�hM��ۀd0��.�k� 2
��e$W@���x\���s�)��!ƙ5\
W�P�PP��w@�_�}��u�D�w�X^�.)

�q�;D(�-�x�P�k��;}���U���:�@72�0g�8��W(<𗷷O�Y��j= �����E�Sr�+��+�`&�X3��в6Ϭ�q##w��._�ׯ�1�5�\�l߾�X�}�}��������z�{߫�$���]:�)|���_����2c�\��.Es�<����#΀�����rs_S���+*��*R�DP=���o�3���!�U=Sv�L
�&!C���.��~_xѥ�?{oe�Y��>{�]c�IwzHw愐�aPX��̹�8� 
.��\NG�\t)2xQ��W�H!!�$9@�H��t:���w՞��{����U{铳���*յ�7��3��ɮ|���A��� ��l� )����[�����1 �!���x��b��w��k<��M7ڵ�^�X �!�.��m=��-��up�+;�R8;&���%l��Ш�w�;x���-��m�52���aOeSfIZ
�Єc�^�ȩ�6ŋELD�DL�	��]�G�2AYeo��@�*u�T���!b�F���k��*Z�&5�Q(c��)s���i�e3�B*u����F��Ԥ��9�R��Ɲ2���'ռRf�k�~r-��2?�f������v�s.�|;c^Fs��9J���9i:�j��y^��C���G��7�ךA��מ�y%�s�yf���J��9��V��V�c繶�����x��h1oذ��M@�*A��_� ��mp�$�~�sx��\?�?kn\)U\�'������>�r���V�6�\u��$�YPD�	A�B���W9ae�4�O|�U��^�:_L�߳I�� K��ˎ��O�Uw�Z �� ���čMQ
l F�{[>��NMuY�)m����("�
����~"��k��Y���MoT-�)������W�kP�y�G��|�jhb\O��y��R�M~�7�c=T25Ʋod��
�@(�c(�bl<���I���¡�Oe`�!a� �&��0~1.�Ȼ� �^x��)�)�nP�}�	s���'1<1/�m�w+�5�)H4_�#�d
�;��(_�y!g��@���wx��pN�A�λ��]av�����	�2�hS��iw	x+���,�76�s�O�B��u��(M�g�p?4a!H�W\�_G��6m,۶�[�λ��3�mb���pѿ���v�|�8�,*��}���
��b��O�?����ߞv�Ev�3��o���i �$p#M�N>S�3bʂy����ӟ��8t�v���O��o��661ލ��s�p]\���z�T�{eh�U���n��׵��J��C����an1��.�A��.˒b=E�������!'B������pec���k^�':hD����P�5�%�=ER .��'�t!|��_��\�/|�δ�u�J =/{@8�t nDm8��Ĉ�׿�-�})���H��`116���B.?)�?��Ow�������b����"��\!"������'?��o}kW�L5+�M���LEH2�d^ٷ�SjӀ��¼0.��QB}���|����Ks�&��<�&�Q�{�~{��;7�fZQvdHs^g���N��K�p�g'�F)H�Յ�Y8#�S ��d����ǆ�ne��h�n �L��?�|�㡞�x�A0_���&��0¼G���ёh����u_�[o��g�$ʜt-�������������:D��<�h�>_Z������i�س�������wo���ZR�zh���V�~a�F��DȦ�T��ɒ��*t�<]h�v�i�>j{�;<;�\` ��o6�G��=�K��@t�Z��7�Ϋ^�*�w���*�A�%*VyOȑ�F�Ď�Di�H&���qe�� e��3�xS���D8D���!��nਬixaF)E�*ڗ{!���Y�� �C��<�@�#y����(�����B��W�W6\){?�a0A$<${"��#80؊~���=E�A�T?��O�{��^+^bh4�94	4��%�u����&�>�\�T��h�t\C�*����&AP&�ά�C�e>髊�@�`����s��΀�?5d����<}�ޙ[�瓋i�����?������v�3.�y��.4�hƌ���Z��f�_tG�۲�ϱw؇w�xR>��}�s͓���P�%�{�� �� ��D���N�CoP��Nx���uVe��$jB5�i^uhI�i����\��o~�C�!<"F��H�z���F�պ�a(�i���6?;e����>RN�P�s��	�-d?�������AܐH���7T#��T`	6>Ă�90�*ϒ������U$Z�	� ����1�)�"���4���B��Y9�"�����
Q�@s?��ϐ�d���B��{�~q�G?�Qυ�Drg��P�����{��!�H��)��!
��9��ClIj�X�]���ų��r�i�ar�9a�`�h*F������u��z��_�-	��2Ϭ�`42�0P�
q���_�����m�Ͽ��?��cR��kVwn"X�f��:�<�X�AVd��\J�� �V�y�~T���ce]�3�XWi�eQ�W='�j4f՛��꙱9���A��d�	O�����R��O\������K��n�9�HNJ6
B�懀�i{SW����������o8����ol
�8
�d8\��9x�"�mi�����7�CL!(%>��!=��#M�BAuVrۈ(wp/s1�:$q"D)�5�ZE�
��D��k<�k���@���* v܏���X_K���a�1	P�;c�Y8@�t�y/����ғ�E�Y5�-�*/2��nC�@�PY2�DK���Nt��%��w40�>c�Bg.y'��0�Y��~�E�+h|��4h^�	L����ݚ=�c i�B��ǟ9r��*�! a���:�C�AY�琺^�h1�s��w��?�A"~�7~�mx0`L��%�F�)�UB{\�����#f����M��'��N�6��I���I�"�r��>O��xD"/I���&U�������~[D�JQ�,�!�mE��J�ǉ|!@v�j���SL�u�!v"�����|�c�C���5%oh�$�8�X�9��Op,��1�*��sH�Ż ���x����,�i]Fb�R5�hD����^������@Ӑ�esк�/��E����|(�KP!��Ar�鏘&���i��^�W~Z�]9�i���
�VQxDI�k��\�c�b��aj�����p=�DJ��h�p%�;��jt��Ԗ��,��)���t"��V7�R��4Qf[*G!�!g�����<���c�a�s�s����5ߩ`#�I��ƽ���L����	O�����_�Q��æ����}`%?�^UL���>Tw�y��*؛^����R沴EO��/mz�p���ik�w\+��7iK����6�s!����Hlh2��2x'x4� |b��$m��8��Gʂ�+H�Z{f��:�`���,-�#y��� ��Wy�@�U�F�T9�0�a�r�4��B�=�R3�m��N0U�15*s/����+*M��҄�H�Q0ϡ��1m��	舾2F�B"%��&,�Q��#/zFz�41d���\l'$G+I]P%�����t�]�fUA`��|م1�O깕/�܈KQ�V�a�SGm<�{ͺӲ~������u�7��.ɽ���ޑ&�%��`��~�<	�Cc�ӂ>��M	�FZ�[�Q*,�?�'in������{��S�L�Üb��Z�Z�Y����\�����,I��z��m��Al�&g�!�gO��A=B�a��*C��(�=i��w|b�_ �0v�[��C��MQ��H�u!L�7��	B
T!�q��v �0R����4 ��3�:����-oY��h��5���g]B�W����p�.A��	��W�
�]�H� <����?�o��R!-b�3`���	�]f��[����L���O^6��Qqi�3��G�G�W��H?�%#��ɟ�I�����Ea_�y@;0,���3704�R�I�)�6k�=r�H�����^���ʠ�}W�����ϼ}�|�~L$K���=�ަɧ�v�yOw?�b88D�+�]f��	wj�s�6��g�䉖2�4��v�g_�m��i�^z���lP;y�}D��AF�?����L���I�-�0�I���I��,����{�����'�r!��C9�9\(���������S���6���0xB�t�E�$�*��?R5s�����+�} �G��!�Ҡ$#��H	�4���:4�s���Ic]�w�����>C����T�{�L��ES��N����n�U�A|r[Mm!*��� "#kߤ�f��@' 1�h�N{ы^�D��q��I��Aȶ³���=�D�1��Þ�d�D+�ko��-��&��{���	�j�����[��@`Ew���<����&�sS���]�ў}��8\p[Y{�,Ac���pX���h�Ae<���$�)�Ms/�w}���|�z�t&����N�2��Z�W&�7"��7������2���#�
j���1K*����q�/����>w�ҍ���f�o����򐧞&�9��呲5���a��ݞ�-�Qbu��d�4����aʁ���W�b+�'��0�Bd��!���NW�p�ͼc V&�:��Ƚ�T���+!�+	i2��M�7i6��& �5/{ُ{��/�K����9��D"f�䨨bދwRn����e<���K;����L���@��y�ޘc4i�t�w7�|��^S�"K�Y�xўpYe� ��V�P�n�&��Ǳ��C��N6��7�4�3� zu(��EQ�S�KEzt&5\�.��pv��m��aۅ1���^j�X"-ƥr�:W4i`��#���8�,� �A�R�u(!�xSc���_�i&E�=����OїZ���Ķ���V-,8,�CN+���?0�v���61J����*����r6[mXeh�#=Z0W��!�O����$:`y~�w�c+��%ɚ�a
@H��4���"�\)8x� �@���K��O���k�%sL ���X��r��; �MP��e��zJJG��i gA�!���`H�e�8;Fd�A�af�*��@3>�x�≫!^&bN41<s�ԯ�q�T�L�H�H�w��6�w@r0!k���f�5<�5��9Zo���-�
�G�O*��N��bVr�;��/ =@¿��!��5�U��Ԑ`���eƤoT͚<r��AraU�G���i�9?7��[�5�Z$���,��&�E6&�����71��Z��KsHQ1�Ԁ�w�N��\�4��Eӄ��Uׁ�MU���׏B��Y�$�b�z0@��B��b�i���F�-�t�fl�+y5k$�����m���?$��Mws�C��P�š�<����Y��Ɔ����Dh	U�H�X�6Ұ\;S��á�� �a�PA&��5�\�/��H�&pp�Va�;��&� =�@�C�\!Ykp��q��t	؂a �cc W�p���
��3n ps�*��H����0R/'EKRO��@����(݅��T:�9H�0 4$�|��(���YW���,�3<�����K��K]�����ye�06�S��-�CVnm���eײ����92� ��w�C�D@��`E�Z���4�V�Z�l4�*�B-V�Z{7��%�C���=)�]�iHJn(�Q���b� }���L{�@/�?��̘����B#]2�I�,$?lj����	��V�d
o�A`+5A� $�B�� �Ky��c���������I/a�h0B�ɓ��Q�j�l���p!��Ea੯�a4�t�Cͼ@�8�B�P1�H�|�DL��%�mAϒ7�pr��J���c�C���5���x�,$y�m��)���˚DF��cj���H�z ��a,<�Ƹa J�3n�@�8���������9t�'�PAY^���L����B���鏌��v!��k��3֒q�n�
?�Z�y��~��{�\�ϐא�ni����\���{�%�w��J%h;���fg�:׫n�o7��ɝ�';\�nS���$Vp�tzv�Ƃ����Z���H���9̛9��ʜ#����#��,F HL�Zڀ�f�����9�Ym0�r��'�+�<j" *l���o�SŽ9Dlt&�Ŕ���i������jZ��e��C��x�V~F>��}7�a���Lu5�yK|c��#H0�?1iw����34H��`��[��uO%��AG�aH��n8�*�1f�_�-e?_�P�KJ����I�$Bļ*���QZר�[,��3��He��3�+Y�=� �\AT�tǵ��+�>�LM{G��$P�lْ��!�K��Bc~�b�\��()]j�e~蟼E$}
����?0�UQ"�0�sn4.�$� �??����ĝۋ�Z�<����-��� �չ@��묭�,���I�d`rp�f݆��ꗿ2{j_� I�!`�8��k9��R4.Bb3ќ��d�Sռ�`���{f�G�ќ�a���[{��:��I��9�I�b�J�g��CF����F��<0��a���`�fa�	 {���������\�ؖ3և�Ƽ�h����?{�f�7H��M�XS�X�-7���D|�FX�E\�R%;l»M��tjD��|�N��N��4ikj�!M4i�b���I����jj��ׄN�����r��@�"�)!@Wq	�%���(��Ɯ�A��T�L=���IS4{R(?\#_��&�K�&C�[���	�2�,ͷ�M*!��6�[g��M�[�k[��0ng���:�����nrJ��sh8F�N!�=���oe��,�FsL��/�˺p���4ڏ�'R�'�'"��aR���h\��	D�'Xyuq+����˳D���W��Ը(i^�&��Y8�dAA��K���z�-h����>6���06�,��Fk�I��(mR�4Y�]<I�������֞�&	P�H�B�V1K_O�C?MN&)[D��P����B���AjH�O�����.��#@�Z�`�(I_k/��ԅ/��Dr"�i!�t�(�X�g���'iB��S��i��ԦEK������(���X��7�nh.��Rv1}���GK���k �Sg�]����:�ߞ�����/LZ����({-_�.�HZ��3����u�x �/�F|y&���H�hz|Ƴ��F�?��/�$ոE�?|MB��v�����9i�8jRW�I_����_���S�/�ik���[�x��a��3��2�B��B��$���.�"�"_�^WO=�	R�߮�g��`v�У�n�X.��P;�G0~�ż�f����Ŋ{3t�����7�I+��+C�6t��_�Մ��`��萪�ZJ�0��'�OR���Ii),�Fh�����Z ��/%������Hת����;D�b�2슩H��~�@�WذRM�=o�j�� &�k��X;�W z)Õ�"Mn���z�W�DsǵbLi��U�?��_���q9+�<�y��(N�K6>6n��l��yf$;�����ؖh���B���~���C��Ԙ�6H�b�i�.�#��g�g�|Ye�䩛}�Q�����~d��ضc�×##�~�/<�<7��ц�GiH�l;�?zj���	����\eC��9j�>b���ȑ�~�l��9g���=�<zȞ���|�6m�h�~֕��#�2	i�+Y)e��$ &�jË��0�"�b��9�d\��6�o>p{x���i}>�w�˹�<(� ���&K�6��8��_(/!N��K������P�T�m�<�f�K���a���n
��H5�� �.Hc�Y?-I�i��R�R�MR�$i��\wS5=u�L��Ik��9�qN��pa�?f#�9���I$<��w'�@Fa>���g��51�T�*¥yW_Rƥ>�{-Ո�YZ�MPRz����ƹ��J�.���K]>�V7�g�1K�;�-����5:uZeO��Yϵ�G�λ�2�Xw���C6;��e!�;^��
�B���L-�e�i�]�����3�58�����k����s\�����l�Ęu5[�9j߹�[v��~�֎#�7�ȁ��/�/�؞qųm�:k���b/��푽�����,��k�z�&��)��6W�q�.�;�l>�4��O���A;��>.��/���E
%/�p��\�����䬽����D�MN� �]�4G���#.g���(ˮ����x(8ԑ=l�tf�ds�{��o�|�0���f��E|�>Ҵ���#�b�"Rq��FUե6O�KR��G�<�h�B�4��u��_�/Ҕ\H$(��K��Yi)Ϡ����������R9+�Mڀ$s��&�$+�O�	6⹂I$aӔb��� ���������jIpW�N�R!���|�[����J����y���H̓a[���{ ��%���>i�cr<y��E۹�L��-�Çp}��8��`�4B]C�Ƙf�u���'Б'l$���h��q.0nn�a_��ce��_��b��3�+��qx!ur�l#˷��笿��s�*��>��O�5���o�T�u�u����!܁H	a�ڴ��i�z���s׹��<W8j�I��,�^�L�">��J��2�;���Zm��mނ�����unԍ�����OHvP��E��q��4�4�Ţ��;%)�9�fg�!w5<E��sK0^1=S^Tb<o+2l����;����Ѓ�
ߖd)"L���EA�~ˀ�7.�"����~� �ȷ|�!�#C�+�I�`=1 =���q�$6�+��1>b��3�m��o^��)����>o�L����5������	�AzG���uAӃ%K�h�i��3�3�^"���=��^O�G�A�/A�<Y��|�#]�N��-�N�f?���m��u�ٵ�Lв��/"���f�Uw�}����|N��p>�v����bXp_R�nX�6��V��x}�ݻ�m۟�tr�o
WG�=���5[Hw@ �ݜ1|�(	S�n��'�	~+sd/,Ե�|�E^.!}�=ca��0E}���u�~/�⣶������)��.�E#�	��I�٧��޷z=z��SY�p��ށ��@<�ʔ �CH�^�c=nsS,Y�А�R"���W� I�J�,���u#*�\?xa�Q
!�������1����<�f5�?aZ�/V2��� ��q�He�Nޖ�] i�g{��Q��w=9y�6�=y|�M����]�S@w\�O��د��hIr��@�8q%ozӛ|O����M���<�|i����q�w�=g�����졠���]�r�ssպ>r0��z���n\>s�9�o�#�|�=Y���'��N?�f��2�r���b����8a���I� X�����{��zo
�0(=�`.:v�d�=��!'`"n2���4�}"ps-�0�`�>�'�=��s��.�;$q|�\��绑�MWg!X4�#�+R�W!"���!�6�5sĿS<Y�3��P�]����w��`�0r��
��DF^?�����(jᤂ�dw�yH�Ja�A�O],ӄmJ�,����0��]��.�=�iH��M N�ϞZ��f�����r'eS2�e�9�	:_�e{��R5סCm|�~�Xs���(�C�I�x)�d�3Ns;�Ȱ��FAc��_��bm)��w�w]��z��9���g���Ja�y?ϣ#Ѱ\,��~᷂�d���*u�M�l&'<��bXu�
~hk8E���;��[�}�1�Ot�_����Q�[Bɯ$�B����`?s��h�	:IS</ۂ;��Ç�ك��t��@�5N�8!aa��!%����	���$���6��A�<Wf��8Q�[���-�Ik(��B�?��9��t�P����w�RE��P�,�ʮ�g�k�sY��V��!���Agh\��܋�QV��TZ��#��
��&�,6#��;�+�:��AG�ĖD0�]m���ޘ"�~i\u�J���hrm:m�6l���-��~܎�[Z�C���Zr.Xs��C?��:�m�v���\�p{b;�Y�Z�Y"�������:�>��KS�$�H@Nx�?��oL=�rcn�ȿv�v�8�-��f;H�%O�q�~ѓ��\�ŒQ��@-<��o��ou��J�KCB������!*¥�tzϲ-||�}�����+��E��|���/G/�����5E�Bx�f	6.��K�5��1�L��eRq���H�8��Ԡ)b+)�)H�g �@�!��I�yF*&���i�J�8�gTq$h���;c�u
xR�0�,���H{~Aw�;�Q�
B���֑����P�{i��5�N����6�.��'"?��/��~p����k����Ş����u�ξ�w<���۴%F���!������Ǻ@q�{o>h���{�j׭�����S�8����v�#!)���I����F��w����"J��+��:� ��D8�f��Co�Tq�=w��u�z�>���G�p�d�+��6�7����x�8:fa8~֯[k���7o���K�F�8V�z1�R �հ �� /��W�7>�r���� @`��$aJcL��]s��@1ȋԽkm��VµsΚ�fPU+8���2��-Rz�W(u7��`����FcG�A^;���.An�nƌZL���%Ė�����3]b+��&��|� �fL�l��́�3?s�����/^�,cQ�p
��{��Fڀ$��(\��U ���F7<+'�b������3`>Ur�4({��}��r�o�]NPx?������-��|�=���yO�V.U\3��)e�UlR��m!J���ƥ6Jҭ���3
sj��?��n}d�|~�W�ӳ UR�Qğ�E���i�mvg�����u�L�>:T.����mf�������W�ǟ��Uts	�|;�XȾl���0[A���^v�Ka���?�G����	�kQ�B�휟�)�oF�8j���~�E@U��<M d+�X�y�>ג�� H�l�~�n\�@4��~�Xx_���ᣨr����v�H�}���E�\�A�07u�٣�"0�b&�#�0>4��۶�w���a"S%������{đ��q�wv�k����`��,�0����������x�5�$E��������geQ�%�#��<ii���)��3`vc�+̃&�/5?�J� ��!M��������@a�	w�v�=D���`�����e�4�ǿ!H�!�[���"R�1�A�|�(v�2�p��}�=7*j/�-�	-���H��@���y�!���:���hI�'�e}��7��6�=�-���z�LO�ځ'{�#y��y��a	
��=��0��[�U��<B>4b+���B���x�A�ǎ�5Q�9g���89;r8�yb|�7.�g�{�My,���@_���F2Z���	۾�b����c��[��={
svȃ6{[��<i#|�U�� _�ڇ�Py�]��gن��mnv��ز�n?x�8=0���䙢��u�]yՋ|s�H,"��� j x0đM�	�x��?di1x�Æ������TPM�?}4�&�B=H9��7!D#��0�:!�kæ�c%�l�����@�k�l��aO$��Ę\-��9�Jf��a`���^Z�$ߴ@����:�%��7}�N ���b�� d;�w�G���CCX$� -�F^Z���y䅣��`�ߺ¯��n	����A+��F)�~C(0C@�
�/�q��ay.̅��YCT�O����uF��؉2YMa�J��ܰU��)b�zr-�C���E����>go�h<�a��/�@�U�����!�̟� ���P�<�g�NU�V׎]�b1��|5��#AZ�gsӁ ����
w�Q�+K��o�F�2B�Π;��+�)�N	A(c��p�Q�,F�<���)[�R�P_������oۺ+KwrȎNO�����OJ��9��߲y����/��Ns�$���vXj9��v��܀���5��l�����e��l��.xz؈�@?�X �U���۶�U�}�o�ѱxp�q�-`�&iR
�#i��?b�㏹��(V`p������!�'�?�CA�ǵ4l�|ۍH�Vؼ�J �@���ߍ, ��-w_��yA���ɼra�b����Z�x��H�lP�~`.儗�(�g��"� ����9$�)I�)���T��I�o�&8���AH���3���'��a�;�d�L��W-����@Z�����u�J&�� �E����7@��?��%Mr��~��k��� ��?����!���3�:0��"Θ ^0�MK�씌�uG�e�L�RV3/�a�d+e@U<wU����|�}����"G�ћ�^w�u��[�Rd���0ƶvݨ5֌�qT���[��� ���5�܂s�p>��͠C�3������y�u&��'��[�/����#�$�}���+���Mm�94g��k��=j��DOd�ư��watj8��h+���w��[Bɓm'<�Ԕ7}��	/�@�<O�����>������7�����U��x�Y�����-��@ H8<O�B��<3��g+��"�Lĵl$
�R:�Z���5ힻo�COl��Բf#fW���G����׾�]�<Z�T�20����Ԅq*~�"z�c	BB2�o�)/D7�Ad��H��F�5N��HT�$E��Y*j!��4Kg
�(��pPyh`���� /��#El*�k��͡
d�J����GՉ����>���9hE������"B$d� ��{�k ����_��B����a�XO�-��3�
�u0vy.)/3~��++�F�f��"L�70���Zs��G� 2����'�����=�;��,���y�� �ӷ˯x��>���֊R�ds�A����6;�̈V�W�U+�%y#{��d�>�����^��Z�����l;���W<�r+W
����gO��2���{l��=���;β��0�s66�ƾ��o���E���&�_��I[�:���Zu�֎G�M^�z�i_��F��Q鐺0����x��Ojz)l�@H<�Z�y���`S(=C��G��`q_n�]�u�ɥdU��k������ᾩ���Q�)�V5F4�[��3|�˓��≯�����UP�M�S�����T�����Vau�9)���)���q�D"T�C��	���i?��-��`R���ai��Ռ?����>�p�yS9l���i���^�g�p{�rL��F�V��)g�4D�[j[`�� %K+Ax���)�.Ps���N�����ξD�C���Ʌ�w ��H(������.���<��"s��!ӟ�Tu-���H�vl9h	��%Z�iI�?��ʖpO�3Ʒ��Q�Wݏ>��(�@8K�h�/�>�-�~#��I��<�e��W����0���w��{~���s��;�|�^b� �0g��@|��p>�v�eW��݀A��@?#���/}���_ז�P�����-�S�ֺ�폎�I���l^6�E]l�u��9;K Ҽcmn$�t\��$k>C��lⷿ����t����jc�[���o ���d�%��qVZ$�`�c65��L!+��-0���{0x��y2�h��-���k�Xz���p�qGc3C�f����Z��	���F�����!L���<@`�/�\�t_�B(���hi}U1gɨ�ajt_v�d>�V�z��`��Щ�������ijo�zB ���M�M\X3c��)����x��|x���<����%h�w �5�ɳ?��O!`���{�����+�3�:ׁ�C�!�h�q��ٻhPt��|�рphh�|�f���rb��>���_�^D�	��D�zZ�|����<p�9d��4�ݤ~���.�S�}C�!!��J���0��/p)��$���������|��a����_���-�ܵ��5�����2`Y�J|p�}#st )h5c�1���������h��:����7?_��x�v?��}�߿�v|d43�M��$��O]���N�����	���#	pPq9�GZ��_x���� y�J�ݖ���_�5,"y����A�}r�3�T6���_�MsU��[�!�܀- 	��i$�N��,��=�q8D^:H�H�ܧ���ڇ/djoJ,i�Xq��P�t�P5�����9������,����RJ����
�������b���]���d��F�	?��s�q/*���9���n�!���ј�Ӂ�	��0�o}�[�>��@�T���@$��e�<���<�Ϙ3�@��<%~|��0����m�>���o���<�,T�JB �g��Ә+�=�va\.�7��wF�^��=" բ<�A=H���Ʒ�F��uߧ}�Z��@P�]F�1v��_�_��~����(@�g�g�D}RT��cM����;�~Ͼ��[��`�w�3�y�B�A�~؞x��� ��'��rWЅ���C�?����QJb�:����&�`�>�s���\�&G�T�M��o��$d�H��ˠ�$��H�HLHe
�`��y(+d7�K�0�з�vچM6;w8�;���Tp[>���+�,y�k���^��(�'_~�����W�jw��N'���d�|���$?�Y�zQ��?�;�`��.UJJ�f���V�y?X5�1��H�iV��I+��@0ހ�0��� �!�z�_�NEf��yF��i Ҵ�r&�њ~\���\p7�̃�} n�� 8,NhG��U^�����}�<,���F̃
��{���T��Y�����_Q�i-
e>�[���
�×�I��{�5i�*��r�`�%A^*���%L]X�ny��9��zιچ����ѽ�������-�:.,�m�M�؍??�`�\���GJ�C�Ё!���M8�gl$�RΆ��8 ��R��F.�^�crk�0�'���}Z��s�V�\I��v⛷�!*`�<�l�NW"���A�'��z���| ³�9{�k_c?��{�U�q5�|!��L��Ar�4��ԋc8vQB�{�"�JC�q۸aKP'��X<&9���k�{)Q��د F�=�2��G�w�t8�O��?��/��s����{�<���v?�ֽ�E��?j\~�3��P�E?�B�^�Cب$0Ta0i���A��N{�e9)4�t�s��t�0�2�ʯ?��&��'���^{�΄xv���(+k~���p~������u׸0	��+Ulnf֦'��?�
������;��soz�y���/{�;��5���R�.����4׿`(E��9�ŰR��bR~����Zנ9CH#������,;m'�B�K]S)Y��|�����sA�:g��߸�=|:n(�sO퉖��6 GyF�0Tj�Ԣ(�Ja���c�q���ȜH{!y�sWo��`��sG:Y_�8��u�s�棞\�n#h�=+)�<�*|'<��*��R�ۖ�< ��7�������"�}�tM"@��#��
��:��Kv�X���Ar��q������"щͥ�h@jogѦ�7M!�R� B���1�~�����ʴ	�La�O����Z�]Z�\�
&�'D���P����*�U�&L����	J�z ��|8���Z�x"��5�,�f@���ۉ�	GNSU�,$z�w\f��q�N���;I�����g�����M� ~r7A>9;�{����TԆ�����B�Q��%,��[��'h��k���b��ҡ�\�RB�+t�#M�j�
ԔP�����۹��.�b��9U�}�������mQZY�EF4{���#������w��!�w`�$UEH䝣w,�:64��
�p���t�q������L���=�W�L�`؃>C� ���z`��4ߗ�+0�Ft,FDy�H2^v~���]�ΡZ+7��g�k"�\�;6����3��#��3������F��)"��n<�u�!aT��S6��
b�Y�<0"�C%gx9D^�00
�h>��3�A��Nޖ�ow��T�b�� �i5�iz"����l|�tX�u�+�=yȓK�&��z�U�.$)�Cl��[,��ڮ~�����+p>	i��5���c��=��l/q��V�'�	_`I�;�x�V��p���\}�cӶb�u��!�$�S��S��I��x$�
�Z���_�B����=�Vn2|��+����O��r0s�T��SЄl$�z��?(& R�ŝ�.>�&����&���G}�:�$L|�B�f������O��HS+MAƋ�ϻa x~!$ +��\|��/�4}�7Z� o��峂E<15C4 �ߵ���m���)%J��R1�0̑�#Vܷ�6���6b#k�ݘ�̗��A������Gr�T!�ԾM�4��*���qg���V|�O���\�rZ�4�*�*q������+xBը�3/�(�5MӪ�J�<�n�������=V��
.�P6[��s80(��
̢m�����ʃ��̻K'�+�B$�~M����J�P�Ӡ���ru��M��V�&�=-+)�1~�S�{h�N*wG(�N~i�"����Q�$d��]i!t���1�g�����!�4 ŀ�]� Oa��y���7�_���o�t���N�Ȗĉ���j��ٓ�r�������u�6�E^�q�}�8B[����p�����mG�J��jZ�+x�����m��I�5�-��޶ԋD��K���t>$]��<$$��`���\"�z�H�0Vmn��~�d'�y9:L�8E�0$r��<_I��X��c-��@�d������=���2p��VjE4��DL!�Z.�YZ��\W���ؽG�f����!u�@�U�K_W���Y�HN���i�g0FEz��k��%�IWM>LHbh��0ϐ�41e,=բg4�Z���px�N���x5k��o�38bs�i/��C	E?�H���`m�s�s�+Pp�m�A���~�	R[M;�u\M<q%�+�E�_���(:+O�]>�*�-���I�4a������?���\ j�	+H�5��0��b;��t�d/��uJ��!��k�@��-��iv	P��ޗ������.3M��p�r$"t҆�Ҽ8+51NͯR�^pt�,��ȴ&����LS�5a��GYYaH$$�xs��"%����"�a�J��E_�R�UeA��Q%2�gb'o�jQݞ���A�G$.,���P{?�z0<�H�{)����T�+0����ƂI "Ÿ�|��Śq}�d���=j�� �!w�=�1��l�_����?7�����vq�*cq8#l�\ڌT�M��$�*Ǐ2=�Z�4F`%�*� -ō�v�el�dÕ��$���F���6�U83ӳAI
?��Ē��V�9%]��%b�������@ɾ!C�r�H�#�m#WB�C��[IЋ<md3P�v�B�Xk&�Hާ<@b ����$�9�v�
`�$e��+6D����������j��N�&AFn��ߒh�Å?<b��~g �5'ؕ�׿.�x����]�/_tXO��D��|�U�����,Ы�A{���D����K���^e��TX�=y��'�9�_�è2*|;����(����cc1hfzzƯ��"
u4���`Iz��O	�
�N�`~f��w/���$��m�}��wY�Q'l�V݉?Iܦ��V��(�V��%��2�����?{|V����� �:�҂䛾��%>�)��Y�J�����vi��
^i��C��u_��O����`���=���Dwzf�/xL�.5"�܄uMZ'���=�Y�s�r%�ڹX�qdl�|U�ȉU4��n��,PP,�S���i6cpY������������Ҧݽ��w$/��^ӑD���y�7�Ʃ@�d�	O�;�)�^��C<U���g�s�:�FFǭ�P�#A�{�὞��۾��݅k��H��+zR��P4)yO�Y�������U¦��29{#��byh�3��N7챃�V]h�T�(��V�+���]iW�טSb�B9��k��Ȩz��jO��ǟ}��J7�,I<�j 6��Mw�P���oqfn��5�]��O��aÒg�`��H�7�C&c�����Od�cCn�y�[~���B�]8�k\�)��'�
���ύ����$���B��֬�Ds3s���cl20����ƀ=i���N�d-�2�	?�Ǘ�>
?;�>�xW��S�n�/��]~�v��A���K�/���4��
]����`�dt�_\�E���na�Hl�tNۢ��i[�U\�y�G�N���U����;<56���1�!5�۱�Ѡ����)��j+����S�O�w��%ҔN-O�'���Y�EϋB���Yg���m۶%�Ջ���!��9'�F'0�3�\:<kÕ	�K��+�3�,�w�K�/�}�C��L�#��!�I���{�� ��fi��3�lu�����);K��k�(4;�o���Z����j����)[����� �/��\��>�����]#l�:���h�T)Lz�"��ٺ��ڦ�6xpɸ���|%���7�t�둵��E��"�*�n�N3t���C�BP]�^l&o��ݲѱ���uWu�T�fe��"�?}ih��(<<M� ����+��jA[��O��o�|��%�L�����\��᜔����yخC�q�����G&�����\��0⮝Ĳ���l
�D��Q i�3M]�r�'�}�G�񩐓\}_��W�}dk-�"�E�!��l�zz`L[����rm$©O~�N|�?��@6D{��?a�#�dW��S;�������q�0p�g=�6>����Nد���{��'WA��{��^_�`7�s�N��_�e�5'E .}^�7�@HS���FU-@�Hi6h%*�%����s �'�-�������0���I�"���*F���T�[s����ک֧-c ���O�<V�˓�$\�-x����CONNۚ��6::�I�<-J�-����b��b������zh��>�������)�&�lg��L��5��}s8�s6��}{w{j��{���wv����3�+v�gۛ��3�����T��z����G+���2�F)}̉�m�= �nn�ff��;��O��������;�ܽ�v�=v��/�ˮx�5k��!���h�#�l�$�"������?��/�c`�t#K����]��g���v;p`�x|�MO�Y��iFEIڎ���A��p|i 2<���(�S�	JS��%���}��j����	�G�,d���o�6q��������z�*��@X�٥�=�ʕ1��j�A���Hު�Bb�����E�%����vw��l7�3?�3.����ܛ���%/y��:�L��$�i�����曾���,�p�n��[�v�z���v�}�:u���կy�}�3�q&4T����}�|;yO\���K.��Nߴ)l8q��s�MO��O�6O�7��2f����_��?8m��ɟv�<�iH�7�LyB��_�Wx`�?��?9�ă�҂TA��y�ۋPJ��߅Џ����n#;Ƭ�+[c�aL/<ݦ�o��Ҍg>̼Iq�����2�k-����ׯ_�M�G�ŵQ�g���?ӌ���_m5�S�T[�en�� ���'���ݠ�E[0'�F1�jں��v�E�:�Ǹ[,��-[�Q�
-e�(s]�`�5C,I	��N������&ug?F�׺g��/�T<+מ�C�=���vn����v�Y>�n�_��z�|�]��gYex��=w��w�9��[o?��;�ߖ�eY�� �w�9�������~sP�6�y�������q��yN�`�n���l���<����Co��%������~��=Ϸj��+H8���˗���rVϼ���#�i�U�]��:Y�x��+x7X��Wng���Ă��O���al�K��O����P����D�"����$#li�k=�T;Վ��׿��;��<���h�b.���7�5�ގiN��6��;�!Y��?����:��I����|�����{��p/��~�4�=��kҝ�|�@�����پ}{=�y�w���G\��ʗ�����}Ǩ?w׎3��;�<��;��?�C}� �E�۹ABŐK��G�c�6���[�G�]Dܻ���1�H��qr�?��+|s\p����o��B�F*öo�#�W��'�#��^|O���U2���}���X�QQgG�qQ����;X��X���y<��@L~�B���/��W���7n<� x#�g���t��RGS��ޜ�P�R��Ơ�S�Q�������)���U�:Ћ�NS���R�S��K�'_Fp�U�ߧe(�q=�+`KcS�ԗt܊9�8U4F��\i_���VAy	i���K���{�0�]1��$�-E�g�]o�]_���!M�R<���)�{����x�����FYG�N8�`���-Y��F��~���'7jYs��~ʮ��s����w<�~�g��fP����
��D֭Y�$�y��]�ن��lٲ&m�6_������7�j�-�����i���V�Pz�}c�\�R�tϯ���Ŀo�K0~��o��a��}��y��m[��������n;q!��������o��o��s�d���q�ڵ���N?ɿ��� -Tgڡ#���U2�p�dxdµ�4�9�L�D�Q�����PM�1���o�#��}���چ��tɪeL�)��C_S�_DB�S��X��mpe=��V��-ՙ[��{�oH@EXD��h]I�����ا�`s�*�w
��whR���+�9H�$���`9�+�\I�y�{�1��d��4��]j��zi�)Q!s Ƣ@4�W���[�S�I�и�GR�b�$��3�-%|-�豸�Z�1�l7ݦ�Y۰q��E���	`�;G��ƈ���6]�-����� �R���zd}���&����w�<��mXw�{��fBok.���M/�[ȕ�H�=w�m?��W{��*�Ɲ�w�b�y��v��N�d����XU�K�e�����AL�Ng)��г}�ͫ��!��0���P�|����M7�@�\��?�zB�c[t�l���=67�f��#G��<'���I7�E͉<�}�o�o~����ZǦ��m�HSɑ�BL(F�}�V{�������	�KlzpP��L*��L�k��"h�LQV��T�Y�.�g�E]��p�&���̝b,��k*ً���J��q�͈HZL��k|�Li&iD/M�O�h����x��� A�&02��5��B�T�Q��<VR/�TkH�N��1����7Xn� j@����h��5_Ms���'gё�Dl��}b�<R>SWg��᣶���m<:��5�Ǖ�
�7�%Y��esl,F��x�nإl#�?s����^�B�LL^9�8<S	���Ӏ�����`Lh8DB� p"dAspG'�"Li�R�r�'��e�(lT�c�ר7|qt�I��l��hZ,��TԴ�js�Te���{���[n����]WP���fQ�vO��g-��ZN����:��)T����(�ry��<L̉���� /$�|��y����H��d."N_qW}����Z�n��!���<� $�RB��M	�E8���ko*���I��N��4'��X�����ԝ&RK�r�W�%MC�!e
),���1�=�\��z�l�E�b�������� $'f��	��>����^�֐��]bip��A�RoTAEiiG�=e�;�:M�N~Xiv�V�]5�o���/�|�ݓR�M�W���B��ֽP{܏e���ZexT��4/���+?��#�#�c��9J���p~p�云�1��83�%�R#�Sw�6O1!M
B�u��9.��lxP��'��i�R�#�:b��G\Z����uu1HC�l�m$�[��Vk̅��݃�f�N�L ��}�s~ )��я~ԋt �����A��v�o*6�b��Z�0�9�	kRM)l�E�6O`R��3����,�v����Z���~�C�f!ց������)/�ą��`�}I׸Ѧi-B"����酂t����m��B4Io�1����N�s%�J*�4-b&��S%u����MꛘIJt�0oiM��_f�#�Ҷ`+����]�D�G�$~ER;�'�j 
*�I���<(��>�K学��Ms &�{5#����2�*�Ij[-��\��z\n�|��*�z�o3�?Vm���p���̡D���I�@/�������Jս�0���g��?�^���\;�0w����m:}K���@V����"i�7n8�?ɮ���c���K�4�{�C�	O����(�b�*�/�����a��g���a7���xҬ	� 'ok�֨�C�<b��[�T�3t�Dx��Xt<f��Q��~ac���\:TIWS��h��S��d±�y�c�
�]��6��Q�cY�T�f3��ii���`��}�K_r/ ��W��U����&�w�Pe����J�]�����T�?H��6R���C��ߒ��{H�ZYkŜ+�j�7ˈ*$�H嚛�r3����G�eҤz%��1N�2'1�h���~�.�`���UW]խ��/����uBJ�L�((�)�EED^k'����:i.S��bAz�$5�ߩ�Ͽy�~`��I���٠��-�l�t+�Dx��O�.E���ͯyJgR?��x�N;��	;p�q_?�w�w�%�������1�o}�[. ���o�׽�u��4^i���K/��|��#���5�"��g�T�u�6;�z�ӂ���iB�/��밖-ըV�Nx�?����k�,xp��]jc#�b�G��l�c�mzf���IĂ���Gm���v����!����&�j��w��~�w~� �R6��H[06� ))�F�֢�I�g�B;��KʡO������!��Q�����a�b�v���p����GV�č����
cÞ��s�׀�$127�Œ��\�P��Qaih|ǵ�G��Ԉ��#|]7���o�%�{!xz��J����E?d���r�|=�S�O�+���`v��u��������������g0~��7��>I���h(���d/�� �J|Ιgx�D���%H�h�A�i�,A]���>BK
ӉQ��@�觠4�*R�+���;�Rږ<���է�^�Do��p:��"G���O[����'�l8��k��f3��2�g��U�f\Pr�𑊯K�:���^W�o9�1����Z�?4 #����m����{�Vu�"��g:���6w���5�,�5���k��Bb'>��dtc"!ި��}�s,$��7o��[ny"0���P��DKk���?�.}Ƴl۶���1(P�߯l lr�5�4��<h���җ��Ŕ��2$��C��������=?d�F�8�p�5'���Ӟt�8�� �>�|�x"�M0n�'��D�&����F�ĀM�
��� �,�k9�h<HFƆ&�!๤��`2_�.���H��@8a��%!�-�l��!A���]|�Ů�+�"̞���w뭷v��@�!>0<�R�qE�h�It4�����A�!�`�3sG?��O/��wa8�^�>�����b#���@���x�'�42?ϔ��{��W�H柹�H�x L|Ƽ���\�#&s��A�b��ꓰ�ZJS�N�0w��&I?�S��A�EO��Ko�f���!.j�x��pK-��?g�N�jW\~i83hay�T�ߛ�eU2�ļ����3c2pb4�����e��A�0Rh�'���a��O��w��q�96_mط��M;x�q����Ex��v�%�k��,n�Z�;�;��^O�r<e^Nx�?����G������U��~����g_ye��Sv��ٶg�#{�ə�y��~#\x���áYX�S����1|��_����.���ȒhW6��5�yM�����Յ�-�����;ǼH�R!˴i��G�.�wo���^0�Xp:Q*,"� !�^�
c��"������5�saTC�s��0��I�A��������"9qX�~�p��< ��%X66`'y� ������Յhn�
qހ���?��3gR��ŕ��<�	.��ox�"am �H��ƚ2<��t\��[�������#���1?�@<��y6��y�X��w�ß�e�!в� �0�J+��z����H?���v���B�w�O�k�����ؙDj��Q�`r����=��nl0"����#�´��5�����9F�Zj�Z�	`�3`���;��EO;;G՘��J�8{��N��w�+~�5��.��מ�c&����?��.�ǚ�ߘOՕ�f�\��0`���c����]g�sٱ.���m:�p�+�a��kk�m�����H�n��˩
:��ۊg�N򖺖�0H]_���H
�2T�3w�gO��{�F٨�����t�MN(�"/!#��g>��@��90��]����)L��r�pl�E�ߴ�Pζ����*�@���ߎ�����+�(>$���VaqK��vߧ���o��*t�&O���
�8C��$^��A��;�⁔L�(BdyLAFK�ć�a <��z�R��?���l���BX����ε<��5��v��F��Y#�0DBȻ �Kpu8D���BZG��`\ya<���0��������\3��O�`2�����D��HPP�l*�Ë��H��^�җz?���Aq�����{�0�fO��y.�/���ó���jg^�/�m�� `�E����Fgh��"L��+���6�����Y�����A󥆯kP�6�`tl��ȯ7�\�/ʈ�%{��Tm�V�9?�N8t��Y�.�I^Br��������������~�;cK�N��g�3�v��}��b�]�%g���Z����O���1�+�aܴ�Ȑ=��>����j߻�6{ы^�O��G��9�g�a��c7�tC8��,I� ���w��UY�j��s?�sV��!�*�� ��QX�b�= A}��a�MR�uLK�(����V���A��s��˭��ѱ�OYA�ѹ�)o��֬�����F�5}R>s!� �8Iud����XUm�[Pb�D	�n��B�!��`y�C�3!�H�D'C����P"�qߣ���2�;#�N����!�2�)]8G:r���C��L߸��>�9�&3�0J�DzN��p�Xb���s��	�M�%�^�s�0�7�=�C������ɷ_�s�b�g<���	k�>��^<�x/ϓ��o�2��I�	�b�0��K��cXZA������vػ���;h�A�m Q�2b?���zw��w�c4�GZʾܰ!B{�G�7�}��Ky96�x��}�S��=�G^`�}�U~��:� ��e�Ұ�����/	�Ď19=h�Hē��q��A_��t0٬D����|SOL�q)��٨���Y��h2�	��|��ԧ>�Ź9���/����!X�WR�F[�7�����4f\M�b��P�e��@�[C/�\?Nl�O��6���B�|持��Ƈ�-�1C�������i�E�Q��q�H� �����ġ��sИ7��?�Y;�c�c.!�<�����!yq8a
4�H?�Fy'k!�O~+�C���x��$�2E`ƉF�{H�"��i�f �<�>\{��A���5h��E�1a'A��11�J���0*ր~ ��,	$"<�*#3sGc��H���a ����z a�AE0C��z�C�!�\#{�y&��z3_�����1�^�g���y�1��D�4��=���RD�S����΃�8;�By��]=��X7[� Ͻg?�*_'�L��g�9��=	�O�T���xff�v����n����Ӄ���Y��F�<��Y\�"��flx��t9�?��~߳�D󲯔��=;�+�y���^��9{$��#�_t�i%s�Ң
ד�&F9n���F�!��� �>�tH叾옺x}�vl??�3�67e<t�>�ߋ��ƭ�A>k�"����i-Vي��ϟ ,I���!��������!�G��F�c�:$Y5{��$�#�qCp�	`�=ćk!�ZS�!}�A�a�H��%D�y���_����� �a]Xs�v �:�4�OZ	?@9����!&̌�A�!�"���7Z��A�Ȣ%HC�9���� 0�����|���<m�Ly70�"M�^��k!��+���yd 8�Q%�A��}%+c��,����� ��|�o��~c,�V�j$�Ѱ�ܧ=���4�����4z/ۘe��y���u�].���gنM۬2<�I�b/#�gj��+:=2�| ��q��o��k{�A�!�1��)F�zMI��~�)�`����>�/0�=Q;�d���5������(�,Wm~n�\�s''��t�B��j1���/���
G��� wN��������Un_<��a�(�9_@9����u��D���kn��X��H2T��Ѣ�]�ɦ�v�7﹉���7<,�#�Qp���6z��J�Æ�@@88�D��o���Ɗ��R~��4\;-�.�7wfȔ߹����bǏ�R}����ɯ^��I��=H�rߤ��4�X;�ʡ�����s���> �L��&O��B�e`�/�[�ϣ�a�`��H��	s���p�>6�'����8`H�M��ɘ��O���y�x7��0�`5/�$�����\9�3Ew+e����@�����r>�qu��b���bzs~
���s�-�	����
�w=_�s�G;����ԟ
C��>���0/֗�����U��4'y��Cl�!ڂvkC�[���ͷ;�w;��ʼ�|v;���saP!X$r�,�c�Ĺ��&o�}���R	�$|�vb�W�h�4F�_��_�_��_w�3�� )�.�_wBɁH7��4���6:��B��!�p<���hƒ/e�7�"�|���4�q�����%��0u$�P!6V$b�{�l<gy���&�<宙F��^�S������C� ~��ȍPy��8$qy��7����lt��o���~����l<1�5�
L#�%	�@*��TiO��f>%,C"?�ٲ�X#��wA�h�B#A����G3�Y�xJK�z�4!}��ZZ�����$Qk�5W\�����8�vC[��J{��-�xK���.��ՊkQ.���z�������u2�	�ŹG�VW���cǝ�9C b_)c�������,h%��w�P���S'��-���\�K�nl��|;$�%�˝r����+��.^��|�qCG8�������A--�Ghg��)
Q��7�#p�x�B��</���p�W�Y�%Q��W��8D��`�N&DCɺn��B$0�}�E��d3(7��i~������o�I{�{�c��G����R�$u�ͽ��T���b�NAW���{�*`2��s�/��*	Sp^%�:�|�HV%HS����yz�,W;��
�V`��1�*xP�RF������� $��Rp}�s���� �Zl`�@�D��adozӛ���4��3�O����f��I{�A^\#�V�z¨�c:�2�k��'��	��0V���}���|ݫv5�5'�@����S��BA9�b�.@i�n3Ȝ�3cD�~P�.�!Q�����A]��ix
�ت7�}���2�6�n�DD*�?��So;	��V*��({����B�|'���R�ͥ�\њ5��� ����z�U8$�T�����ẇ�k���~w��˳GH���E6�.�K"�px�T�:b��W��'�nY�`�R�s���L۝�H�TAD��0p{��{�ԩ�5�D�%M��Hʥɏ;M�JҊh)���4�l*zF��&��RI�&��&`CW��O>��VD����oi�`�A��-f��c�g�)��h��]ஊt�D����ް��w�>1=��T�M��2"��U��[�-%���_o�~n��-�)�c[��3�/0�@�9����p����~��ֶ�y��M�f{�c6ng�n3˻&�7�F3��U���� cFg1O�W��񮶃���张̢0E��R��e��CY!�N���2�b!~��V��ϧ�+�\�&��Ri�Z�Z�v.&�r�' ���B&M�,Ҍ�:"N�p�5��:�{�����?l䃇��Ƀ67{ت�S���RD�$��v��5,�)d�I[K���?�%�J��Y`�TAT����q���H�H����C��xC�O�囘� �x�=���E�щܐ�	���&?�7ݣ흤�D��/4lt|��v��*hxl�S:S�	�A��k�-�BSFtN��i�i���\�f@�C����w��#��Q𿛭�f�t�
O�v�$5�jC�Q"m�W��w`�O�V��b��XʱPT*��E�)%y��3('�6-5�*�w9�Qj�l��8���x��c�Xo�@�|� �/dϴ���$��9��)#'������ϵ��q�?��=1�����sI������~���o��0��1�H�T���[;&v˵�-aM�%f�g�=�����5/�a�Uv�}�&�gl�m�7F���kڙF�g�`K5i3�UE���������vF��Eo�J	���\����^�|�[�J���d� $��m��A����S�q@�C�OE�e����� -2��S�JM�y��;���}���{S�}+��V��sso��9�����k���n�bwio�ji�I߽�_�w{��٢!(�8� ���=�y�8�Ѳiy6A�u~�l1���g������ ���o�׎?ꖂ@�y��`o��2"�ԭ�x.\y�%>c�����,b�CS�y���t(�"xMj!�C���� ��$E��ԷS���(9�QMk4�b��?�JX(��F�.��U�U�<���^z1w�d7�HǆJq�w2H�c%k4���)�.#F���2{_5�q�8/�Kl��٠�F�c.�[�,�1�[��[¿���{r��{��l��7��1�胱��-���/|ZU�jH(*-3m�F��m.mBY|��ִ�����1���w���ش���5t2W�mgƎ>�@�1����x9W��C���p�F(���K=�۟�7��(J���=J�
�5��}�m����(�!C���H��t�8��B�^o��C�l�S'-�rm��6��=�l߁63�g:�X��ke���BZMk���a�-�6�e�f .5�[/W0���؍��>�Ϊ�1KY\����l��_w��h�:��V ��*^� �8b���.*}�LF
��C0��'UX�s�=ç9㔰P:C�i6\�ѩ�C���J���{�z7kh��K�t�ދGB��&�W �e#^�R)2��Gy�i@��c����<��o?RlyY)=�S)������x��V��xtσ֜���Y��#�{�68�4
��c�`��h��9�i4�jQ�ˣO��c���֑bX� L�3zx�B.�(���p]O��f�GP�L���)�8��ӛ���pH�Y J�І���u��q�6z����\8��H���=���<?o�*�k���$ɷF�:ַ��M�ۻ�����gN�sAX�mf�4�jA1�4(1}l��u��l���^<i�A�GDe��l�m��Yrɹ��+��t�b���S��!�I+!AB_�~���X�ݳx84ۊEu#�a�U�ޖ��.x4b��ʵv�78�?¿X�� \�ctXO]�fpl�Zq����e@�H?�W�ݣC�v����ڵ��l	�DؿȔ}���:~���QF��l)�xQf�g���w�7;�9�(���[��thb����@��P/FF�o�s���դ)r��W�RC�9�R`J�y�K�q���_�u�Ycf2X'eg�t�C�+�q߾�v��;���	+v+1w8�~�3T0Js�(FEX�mW�
������� T{0;?��� d�H��9)��;;��-�'Y�m��Mv�5��=��a�y�aC�5�޼�;�o�s]O�hw��ʷ��O��Wz-P�����W��I��~R�N�_��_w&�^�9�?ˮ��*۲ꐚW ǽ�p���;wy<�{��.���ډ3�+v���x<��z�>e��,�x���꫟f/�����#�7�b��N?A�5:u�t�F��M�(`-$ �!%�L 	w^G�� �����5���^¿ ^9i���A.�?iǚs*!�m,�ȩ��SA���S�D ���}���g
R������?�`8C�sJ�¡��-���6�*�v-�5�d�<=���`��V�����1���E?�9�I�����2kU8_��ʏ����W��X%��9n�	�Xj��߲ҕ���	�ѽWE�O1(UO�ޫHOך>�����T��Y=c���2�^�:lB/�b9X�e
9�� h�M�c�a�XS�x�b"����V���&$=��/���e=c����y���ʯ��i�c��q{�w�]�4z.�����0�i/Ɯ����aՒ]v�v�,�`�o�����OkI�EO�%�Y/��/K��i5���`�o��K^�"p"�v{����o���M���~����.��R[�f�5�mgy�RH�*Q� �P<7}�o�[�3h���^+�����"^�q�	�L}&,Jf�y��۴����=웶������8
����t���Z6"H�� ��Vo�TA�f�k�8m�"�Q	c�$�T���u�W�Jx��ƙ/sRe�)ǉy�Ŝo�!���L\Li1��sD�s�񚠕4Q@<>\�^^�x~�)#Jկ���� .C�E��1�7�4����ž��(w��n�����7��Iqn4fmr�v�jC��-Y
mv;�,ve�k�f�s�&����f�n�F�4�������3�8�c�%;�԰��:���S'�ѕg
/���p���k�pf ք�si"��9j�zw(w�;lF�ú5k�&��z���Лv����W�h���u;~���DXl�w�];�ˮ�:�k79.�u�۱#G�?!�b�r
7^���|�+_��n}�m�h�������Nu,���!�=��]�a������lf�D�\:��6���OeHx���={���g��>�����݅�;�����pg���V���n�
ȕ�W�]��x*P�P`��<��g>�Y'�b�_��BO5U{C�!�̙�1�&('x:<g�X�����wZaxpD�FM�g��5r\|膁渖ok����"(�����4u1?Xo�������q쑱Q_�:?���D��A��uk�z�0�����gW@w���p�T�)�߅bֱ������ׂY�z�:[�bC�#I���Q	�:��kϟCDn��0��a�Řbm.J+�e�8��m���{���ҿ��;��!U�q�5��u7��T3�^z�S~�C��1�J)M 9��_잣�O/˟��Y*XU͸�ᡟ�:IbU�����^5j�.X�<:�z���C��׾����v���C��!��WJ��>��hr�0<(�U~�'^�^	���C_�<X)�ël��~��{�}v8,".��N�F���cq�g��i� Z�<6@���kEB��B�@���?��@3 m3��=z�K^����@�c5!�9��P(T,u���a� ��)�a�y9���պPMVd53W�)�!_�� �Ie�o���qm(+<<8͕ J��v���p��;�A^m���C`p?FǆGFI��������X�Pf����7����\8�ڱm�Si0w�k��͚R��<�_o)*��d�cࣣ+m3m��(�f���n,�,,��0$`�Ϭ���W�Q$cH-�'���>�g�� 2����e�U�ׯ%<�o�sή��
��w%�F���O}�� .��i��o{5��?���v���7����/�3X�q��:��YK��_����Um�u�o�� �&�R�88¦:v�MN�� k��M.��x����8�#*`�QYs����y
Xt�z)��u����EpO���-�u� XA?p��V0���52~���;|�#��H�r���2E��X�m'����~�y�#>���ѹO|���� ����[�l��,�Ga �x&��s%���h��q�5kW9$ǳ�y�]~�����\�q|^Ûcsc��9#����(����!���k�E����-QT\J��̱yM� mjR�|)�n��5ǽC�n���Y?NW�.��Șٱj��{	�V����q7��m��I�J��P ���{�)T9P��s^�a�7rl�F
=��]�z��q�����=��ɣ��r1��k�s�3M/���b�䄑X���������.��a��+��w�;�����/���gݶekx�-k�j�#��7^ikVӏv�ff��=�`eWmo��4� �og��+M==y�~���E�B~N�K��K�sW��)q�b.�^����j�����>�KG<b1/}��Kv1�VӨ)����'%KU�(�#�Dt&FL�����-�"����/ӿ��Ω"�p���J�yFT�JC4'������;Ne2BQ�Xxfs��~L�;׆���t���N�^���nܜ�&�0�3�=2=x�(
Un�lX�^tA @����}�QkD�+�{3J�/�>;���ZA` ,/<��銻}��6;q�S�[(D"8h���aO��ۥ#v�nŘ�O])��)���;��k�u�4g�A�¡ D��*>�z���Ԥ=��=�rŰ������#���v�G�R*ة'��ذ�B��}op^���z�g� �z�_��Rtv���XN��� �N�,����a�@fV�F.�"��v=h�a���dP#���Q�?��?�M�Pb! U ���Xo��|_��d!(K�x�Ҋ�Ƭ�*0�6�њ���ɰ ໯�p�.gt+,��l�B�yh������]X� e��������X�,�f�����P�\;K� �5&x*J�󲱸'p�K�=���~,0��g~�g\� ��g��fR������[�ͥ�s��=�v��
�d�_6=�k��g�ry���kF�?���v%����'̕��@�̵���kc.bC�U3z��2a]�X�W�s�p>�g��1pϸ/jCyn�QH	tm1�?)�<�X�_u�W ��=yb�V��|��6�L��I�pK=���l,�6/eee1�Y�@|�4s����«{��{l��Ƿ:�g�E�p����S���0�B,���W�<��̉���?�y��IY���(��̔oڑQ6����A*�U,Kl�)��iz�f#�T�u
f~����R��y�b{!��c���9;tp���}oX��66^��k���E��@YZX�۷�#C����+A܁�@F��E���k\/��DM̱���5���N"�k������:΋@�;Vp6��c']�#�Ԝ��،��^����.3s^�zE313�XPףt\^G�)~�@�o�r繂���|��Ԁ럘��������Vf���G�P&x��ȍ�qn�w��^
־�1��	؇�T�8��i�FA�5.͖w�b�;~Ć�ﱡ�UaM�[��{��k�#���S�����
��������a�������7����z`Ȩ��Ӛ���ke�(z�d��"��"�@��b,qxd��Z�"W,O�"���)��>7��l�]]Z'���Ց�)~=��K�r��[��7l��%�V��p[�l\�����?�������\y>wki^���e�?l�sAIET�3g	��E�(�"��ur�[͠h,X����u�0����H�s���j�
V��/pKA�2�
e���~b#x�pB8��`��^�ʯ�?~��杺���[�¬1W�k���.�q������#�jժ�֨ovܡAM�/Ͻ�9. 9��ب7�n4��ޭϸ�ߓ"`�dg���}��ܺ���+"$�7�.Jx��5���O~}ܓ���%�l|�F�m����k,���~�w�r|��Wlz�7���;��B���r�����(��[�9d�<Pd���/�y=�Y�v����� EI\��0/�~AJ[M���<U��0�RC��& Ȱ�qTӡX�֧��i���TťF�!���� �뾐d�p�[����xk{k�T�e��1[��v\r��׃< #���S1hɕ��q�Q�����[�?��'��\د����ۯ�����ҋ/� �����)��JT�%�@���Q�t#�X��t-�W�@3�ylx$�g�T�K���R�y���j�W�!K;���vX��9�k�{�iG�����w�k��9�U5�E����ի^�P�0ؼd!�����j+&�Q!m^64�D���>;z����e�*��$T�˖�B����Y�g(�
�m{��^
 �}bO���0	N ��և4����pN��9�Q�/֋Z�?�wP��,&yBx�2�a�s��fD�'�+X��u|�s����C9��zZ���1����J�L�5悧!aԣ4���f~��c)5��B������.�E2o5@W<F���Ҋ�MxWR�D�K��X��� ,]JR���v��z���PŸ���R�.='N�f@�3�^��sL\����(���8y�{�T��'�Z�S��k�(_������B��~Ϟ=�'�'��׼�[���-o�,Ω&���W=ﱆQԫ׭��bSӳN�7^̮ەV���ȕ�e���Q8ݵ�Ϡ�Wp��b�7��W<88����_���pݵޡ�۞���C�e0n���uހ�߰2<Ԫ�;p̨�A����K��y���wz0\�\v�BXW]s�o~`m�٬� kyfz������f��m��a;9=���iD��r\� y�r!�+�y��~C}dU��o>?���`�"�����`��]�U5C�H�_�zsU>#��&���yO�T`�X��6���P�����>|�M�5�y��F癨Z�g�޳�_躽7l�M�1���|�P��96�������ؐȫ�[V����^�PR�Zi�8	"Yв��B�@SN��	�*ӊg�ȩ��e��U�:w���ɭ~>j�����c����W�Y�4΁�H�H%& v
���DY�z���H�W�4��eu7s��\�X뭬��@'�?��'&��|���.�](؀��2��=i�&gmhxܠsvt!�Y���7���}�+�؁�/��灂�"Y\��H���"�L�.9�Ë}߽��ϼ���Y�x�6����AV��]87���[��E���s��n8>�?b�T{F�Ӽ��O+6�!��bx������+e�ґ�>�屑!۾m��_����:x�<�a����CA��=�U���BV�������.�!m��K/w�W����&vh&\#�3B�F�@{�	��`8/�
�C	�0�xE;Q����3�u)F�2�\�36PP0�	e�<H��~��x<���o|�=���Z�(pu��N �{� g(�����q��|�����/��9��F�=�<o�d�[�� 歴����=���=�뮻|=)�V7K�˛J!��}Rn����LxJI�8��RPEw
󤰍��������+�,a��+���-��!�+� �=X{����_�����a��iZ,�g�'�{�}�^����~�����R%�ͺ-�o���@x���<P��Y�����u�:�sb �Y�x��o��M�k��|l�~�k����4�A�tl�m�y�%���M604hS�s����B����g��_  �f��j���ȋ�O|���[���m�~�w�yd�^۵�A����+H���˞f�_y�]|�����qc�k��h��_�W��y�L��E/z���%
�C8h#�z�ڂ�ynz�>��OZs��!-��1����5@�<������`��]R��+��źP���z�k_���?����� <�������T4 
�J�K"P�%������Cyb�*�&�0L���tL�/�D����gȖa�!Xو(���o��m����i��{,8Rq�\?��?�0X.�h2}ڲ�Q"�x���.8���T�F�=YK(���7��9���7�1���^ )��e��%lH��f@�Eֵ�q�P��iuu<y6�w�
l�C�N���dm��.VZg2���{ �y-���?6e*���ݳ��{����A91��-/_�6+mbr�ceP����;mF�����'�vvO)Q�C��d�Gq���+5`X7�x}�C�֭�b���>��]-W|Τ��_�=�����z�&��a����g��q�q��~�
ݚ o?˹F�>��Ϻ۲��`��ƛnJ�{��~��`�+׬���.�e�"��E� ���ᘈ�������rx��a��Y�A!�$��<��wx�w�=_����`��:�!�(�u>zl6���rh!�Se/n��>�-/�1/��Qn=�M��MДkG���6���Kγ 12�E�	�b3pl�G�V$���*����̅{I�%n/
��3��=�H���B/�����;��fnT�FOf��/ރ�Ұ�����`����VQYH̓�^k�B����O��	b�S��Ҩ�F��'� ������[ǂ�u,>�='�h�S���1�*W	qF��W,@�[�B0����Q�<C�-o�����[���ӟc��1[�r؊����ʞ�I�;�=�5�6���yn��K�o�} yld��R*�'�w�?\�!��M�X^ׅ����FQ�$���Xx��֯�U�/��n��[w��?u��2��o��6m���0�w���ѻ?����+�Y/��ֻ�;�T1p��`�~d��ٟ��^��Av���k�k���HŬ�:��X�ln�VA$
�)��`RV�\������tK�E��������w(
B����Y�Oz��T�f.;,�/��S�V_�e1  ��IDAT�9�N[ذ�������
��=��3�&�
��,|\�T����@�\#�8��1Ҥl�(�
!���Ȇ�ް�8BOE���Gys��e�f�R�����h�3�g��E�rI1rY�\�,e:�����~l��!�Y#|��B��s=��ǣ��Ul�$DdK(J Kp��K(+� ����
�+���4{DB\i��e����|����$#�y�K橸�2�4o�)-EvU���n�Ev��WS�y��V���gf���[��+lj���1�|h�X��O*���tO=#�򛜎�is�>g�췗������~��z�Z^EVpr�{�����^��^�5<�<X�+l�E�mnfֳ�FG��.�+~�#=�ȁJ����9w�8v{��O����N�� C@��Y��@,�w������n��6�,V�ɐi�,��Y��>v�G\`i��0��@����q���Y��=�x�;��X��%J�%1#E5(�JǙ;K���
E�}
��_��]gb�D��oȃA�2#�	sF���#\�����pl�9� �V�ŀ�&�{bGDx��;���?`"e�7/�����: ��6B�\z} JE�[�����r~�q)���
��X��^��;�c.̕�t���qߠd�C�,��3PSp���|��ZB9W�U�Pe�p-|�����P�fjy���R8U��"0�#�B� ��#��*��uy|(��� ���y���k�xf\� ��?�A���c����8Ć���}�T����U�"��{h�f�Vۋ�ʵj�������E��@V�u(F���5�������]D�X�y�S�[����g]��-��]���62dM0̠�����=�v��G?l����3�ckiI����6��ހ0�&�ed�<�QK����}&XjP ಣP�G�G�Gz8,��f'���k�"E� ��q6�d� (X<��ۿ���i^�R4�u]YMMUm��	+���κ���wߧ��r�c}���c�C�{���@8^x�_��}�V�QH�D��9�"�6 �S6,��������TF�
������
G�1�!����B �>�dc"�`׽��r.�P%�|�7�e����>��7��
�p�@ �!�U�P�?�˵s������b`�PM0W��'k=%����d�=��FW�X�y��,U/�kn��V��ز ���Ǽ喙0�geYO���{)���=��e8ʑs��Pp
��.�4뽖Ѧ��R������_p��l����ɪ����2͍���)��[#��s��ǗŶ�@��Ś�B�}S0&/��J�X�������͠+ŮD�r��q�����,�L7���k����` pe�{�.?PQ�9�5 ^Љ�]j���
��?�!�{��͌�˩�x��	�]�ͷ4,��dq��45�ZeC�`�������/����O��
,�3�����Mn�⡽�>,�^�V+�>��.w���-.��5d5���E�@pE���:x�+_��닻�)k��]@����`T������T����l~��jV̣��:J���	kW�+c�%��W��7�r�����ͼ��:O5D�U�&�e{`щ���'�'�G��֑��T�(�+����\���&����J�w�f�Q���hrr�_S�XP�j�Ny�"!�'�|��"x]�(3k���W�*2���L��u�
��B��_R؉������kG	����5����J��u�&[�vC�C���F�f��2Z�ڡ����=�p�IH�0եp�����T�Ǌ��=���S�>�;*ume�Vx
"����no̿�]�'�]�5�e��Q24�7>ZT��B:5�� �X>���M�<��M�Wit���k��`�u�b�F�����Nc�n����pz:����H�Q�
T
���B~��2L�`����� ,��?P,@-Ef�Nf�7i����g�0r�<�ShcJ��hKA;s�ֲ�����"!��+y��z������*|�^H8����dR�^�J�F���q}�#c�-%����*^W� �3�,87�e��=��o{�E2�����`�c�
�K��p������\熍�eW\�ﱽ��t���=�����u�����f)�<�/$,��"�U��i��vs>�薧}�+
�#�?I���_z�Vw�����g�#>\��Aq�U��ǟW�]�٨��+k�_?���Ŝ��=�=8������xj���6gJ�Y/����q�t�eeҼ��n{�MۚO�K����nXWX���z˒����K�Y
��z&+����)g�B��Uv`��� )�>�8�AX0X&���gr\�,P M�N,<�U���lp,HÁ8��9��8J`#ă/���p��b�*$��=T�
�HlŋUJ��x��z���,�� ��9�I<�(���x�9�+׎@d���/!�g�G���cP2 �Rذ�|�����ٟn���z3��7� W�UB!�V��WU��2uXlz�9�Ph����
v#��\|����s.����꠆ף �<�����j�9ǥ�u%��5_���+��ݏů�n�#��9�ei�Sa�<��=�z�Iߠ{h4;q��b@5镲 ��t���)���?�'�5�<P*ts�گ��BLKu�"�X��sc������_�a�g�-�j>�E̕@K$K����<�����))��=<,R9��~�^���yF�K��#�û�M-gF�5�"��W���^2��,�Y�W�&��{�U׸ %�K�
��I�;���{�\���Gq�7	���0J�+��Pmx����;��L}�
����h��LP4�B���rl�N)�B��CJ�� ��9�
����5��X�j�5�f�w������,���

�`�ū̚�j5� ����x���� +J���2�!��0�W������7����1�N!�̑�@�F�P�iL(BYJ�-o.b�B�F%��'���y�*�z�b&��B���S
�̯����ql���(ԭ�l)�<���B���VF���4+�LZh���U���`�n�/�p��m��gPP����c�I9) �,��^@�s�e�� �2x�E�����F����������p.\�au<_�=���l�ѱ�3x�:E6E�S������M�/]kl�"��d��ĺEp��!���۵k����w |�4W�늴J,o�K�t	*	8��c����y+�4B����_A��H�D��u��7��F�� w�X�j��2R�s�-�5s�(3���ÛA90v*��!�D_�y�����+~e�(@�5�I��$P|�&�7����hE�Y*�|xA�?���\��E��d��� �h�����Y����\}��2���,.%υg�ץ���'��f��ĜQ�<_M
�i��"�no/6�]=����Bs�p�C��U[�:�̍���9O���Պ�n�� �<G}L����5������T�d���h:��E���0�b�9Z���?�������9��3Y8< ϭ.ƻ�ng<&����Sˀ�|`2D�'#b3w��  �c�%�=�J�;q���}Ȏ���
V!V6OS��-�O'��S�TQ*X �4�a����Z�H�!@����4]EFlz�� .}>�1�TʒM�<��s?e2�F�qQ8X�X� U_^��\�x�;�ax��L
#�J-�\��5�=�X�y`=��B��� �a>QAY�YLɬ vz�h�z�:Jc�+u%���c�O��&��5 'I!��<A�xR�>���m�>�_1Y�xO�o�פ�Vz��I�H��!�J=���N^���w~�b�b[�Jl{X�1��	*����.�r�_#�V#��Y+-��n�'U���Ih����x@�qnJՍ��R��]�օ�g":����3�.�g���������6`NY�-��}ou������W�7��).o_�5�$ L���m��p
k����c�lr☍��j�#�2�}��+͔�gyZ�!��<�����o�'m���%s�_�`�>��Kإ�����"l��:�G>x@-�!�!�KU���e��"�
���!��+���%��2��`05������ �X����=�n]*fJy��kd�xR^�zRПav����L��!��)K���K��Q��k(t�T����������ͣ�"�w���3n�նl�(�����~�a]�ךd.ɂ-'�l)*��g��]����������9���٨ (ҀX�N��)���nVx�S;Ik�">ǉ��{[��	߲��4��h�W$ռ�Q�h�~�w�x�2:a^�v�;�6�E��_7�s�ȫ7��r2��S4[u��|�U�q����NA�,�>���i��$�ѣlwb�03�T��5����A,���p^]y�l"��XlY}���V�v��c��J){Eo!,�f�b���=��٘�e���@�|A#�a�#���������6� �p=�{ѵ�]V
!&]τ�c}�#OP% FL= ��e ����Е)�Fձh��|�ǀ@�~S? U��ൠ����|AF���I� �@m�><M���L�Ac��&hG�>ץ�]�,�@x��s��f�(0�BF��f)\���0�fI	��N��Z�����ܴ�����~�ɩS.\f��5W*�zZ\�
p]k��n��sn���W��� H=)6�Ou�4%��$:����t�3���m;?W̕+�
��O���^~���-W�P%�ً��'B
u����=/�?35�ߋf���������-��{����F*��-pE�9wP&���t�)���9�X���x}��۹<
���k9�D������4#L.ndi�ܞ�8�F�"��z-���*���)>����^B?��+=u=a=zd"X�E��� h�5�A67\�z��Y(s��7�6�(��SgScR��,0	8��.X��M������0{捀U����P�g�����d���je� ���̊���s`�@7���~���>�<��96��<,w	@��T�)m����A�)�ϛ���R�����86�'�+�WZ�80��ԪR9�R�R��$,w\�.*�ytM�:��w���o�-�̇�������yC�c)���3�"D�\�=�}��
�����kIXCs����y�
r�6@���	�[z�L��,jf6x/��%��9/جt�г٘�}�w�Z����>׾��1sϫ���(dJv�R��f����7F�e�s��'O�c���#p���-,h��N	�c��Z�:�?����oΝ��;W����nӘ��3\���2F�%�.h��\�^5k�*?l�Us>t����e' א�'�[A1Ǣ�D��t�?�͖��x��a�
�xF�\*����U6[��M����d����[x��s��s!��p�4��5��'Rl�G*]/~�	�� �W.�R�<�e�I��}��bl�����	���X��A�my���,�f��EX����+�y�0�����S�B�_P����B']_��jϿ����#s/4[+��S�H�&��p&q��<#�%�;�����{�>	x���(���Δ���bAZ��պ��y;�W�$u��IኧI�N�������&[����{eͶ���q���M���N�\��{-(�L�1�b�i�펧���?<<j/{ɋ=A ��b^�������9J��^�g+�@c@"W)Ÿ��̔{Jp�7W� �9o�ĺ���q��Ɏ�_��������j�@�}����y�V�:d�@�w���BD
,|Y<
���O�X�T����,#B�-�������Q;z���;�E,�V3α)�FƖ�l�aC���A��#�U��֏Z��+g�4�X�??�@6�|^�b?�-A.�T�\�Y��LBL�.���\��#!�znj|�"2e�nR�+��\%����ϊHB_�A�H��o	���ы����(��*�!~bg�Nn�ׯ3:����J��/IC�&	e�-`.>����{)/����o�)����Z�B�����C«�d6q^���`z&�D�.�
G�NJM�a^��V�z�s���a��lnf�s����䐞��[6�Үw>���g�
8Oɔ��o�s��L��=�g؋^�b{�[���.�w���5���ZԞQЛ�B�əY?���k���$��Q��r�a�}�p��Y�7�Yz���P��*@���ew�U�r�j�`�\*n��_�����S�G��6��Y��cA�o	Yy(8����`�B�~�{�ч�e0����Y�B��g��{��y�a���K���w=#������x��k .Y^�Aۮs�p�'ON���H�јuET(�l�ju �{�s�*�X���l����`���BX,�
�!��Ț!HŻ�e0J����}�;((6��Ș����ȣG�g��M��S��>�h���e������ �v>����j�=�� �)z�(ޗ!�w9���k���0T`W0�`��������e M��DU8���9��;#��s��/���ۻ�ֆ�T��D�c�i�P�C��p��GF�TfAn����3J���V��@,�����n���Ea���Zv�����M�=�r������}ͮw�r��(��|o�˷9��1Q�P�P�� /�����(C��L�FO(���O:/��7���8
��# �Y�G���|���E1{	:���3��H�8G{�v�0$(����Lx#t�կr��a�V9��Lh�Ć��sa��'�&lU֭�>YK��L)�rs, �@�.)�i�2��j����@�.��V�;l��I���]1��`�ݒ�x��>+@�L���K.��5(���ov�"�2H�)��9�k+%S|/d�|�w=��X7��ʓ�(�����$%��$0xj��UK��%?�E�%@�(YJl.��$��&'<o�2!���,|^�:���%e �;�Y�E��?�"��^�qI]�>�*��<H�Խ��|��� �h,t�di�����}�(��	]�&�&����1��{��E�0_�����U����K+Wr1���mr_�kN3�� �'*ϰV�\�$�/������^h��2������9gqu�C���(���LLĊhkG�\����K�-˖۝/{�C��aR��c]��e[�f��ر�>����������A�]��ȓg���7�ǣ�x��٫^���za�fc�EK~ �~tt�Ɨ��-�0�*h)��1ɒa����E"�EJ0T<X�l`�}ua�9=.���W�,�bݩ��S,�4����\}*K�+�5C;�6��aS�ؘ󕅧�m��s��J[��2�2��AKZ%�A��M�~�(ā��E`Rp%:,Yb(A,"�K�'J!M@�cq.�T�у���TL�� �Q�(-�[j.�0`ŒWz(���Qr=	�r�Xn;�����,f��=�؍�B1�bD0���W�<�j�@��z�����
e�\"�	�4՘!�ε��P�j�.��X�֋��GZ4���j�Y����/��/�ڱ����x���;�d��������f��1���Pg��;'�,�P
JmOi6��4��i�}�I�+*��h�N۝�M5:��S�s}���� 2SN�Y�O�Ӏ��oϞ��>f�)���W����ړ�K�-�hX�ϸ�&�pi�hjjjL*/,c��j��9�U�8���)oϪ��Of���!�E�f�*�>Y�j�����{Ͻ���v�����Y	s%<��o����&o�c�E�1�"����&��g�gsܛ�A
".$.6��Rz�F��U���r��E]O#]�|u��5fO:��C>�*yJ�Sp׶P�Խ��W!��(�兒�|���UW�k���9#�j,N&V1����w�6%��M"J�h=E�%��EѢ8�.
��x��PЏ���pN	p6$B%�����h��$� ��s�������>���{'��MLsn��(R>U��w�f��1�dF�b�z?�M��:@��ޑ�z���2\R�����Q TEE��S�Y���KR�1��3KV�iv�Y�C�K��7J�NuY�:��KMg0�����H�����'ҘA�{�&&�����%S��$��
{�ہ�o���.'W�+|��J���
t�{�A��zXC����x���opo�����"��P��g�S�K���v��kS����#�/���o�kxN9Lz�u�������{1zX���G2���n��}��;ۇ����A�_v��v��O3x�[A�۳���_m��a۸�r�T���%���gϼ�v��W��@`�R8��J��(��Y lr�����l����-�4�s��-($kl��m�z�f��>n���¼���:O��w=��sY������a(���a�b�"���" �0X�@���{jW�k�@�3 -�{�E� ĺ>�7�e���`�J�?c�ca�T�~���Y���&eǨ��������� #��|�NA+\�j�9�h�sǺOy]t�P�<s ��84\B^V"
����?��� ���	�WN����ZZ���k�Z�>(k��9?���Ȩ��f1��S�ǳz��_�`���ՙN1
]�e/��4;Ią�����1�`���}���U[j��>Z���(���6ۚ���_a����C#nu:��V�I�����E��� ��w|��W�Ws
�=q��N[�ض��v�׾���
�t]�+"�i�БÏ����{�9w|��_����M7�b��~�ב`�T������/�����ٺ����M=����o�@�����8h�.wpjj�N��6�χ>�A�x�� A��sYQ�Q����	k���X�i%c�٢�z���b� ��Ҵ�e�e�k�7��2�x��0��sb���u��ӿ���֪Rf����Y����9?�!�U�L,{�9���_��s�4V5�� �ʔ��ō%����gs!D(�����a�X��<���]'X����y!��c�i����!��(&��uE�9�r�y�¶96�F��>����R��+HY7�(�aH�������7bJ��!�eaQ2�0Pe�}�e��:���a�k6����&\��;����2���dw���\�,y"��bAٙ�Ӫ�Փ^
���\;�|ݰ��s-��+�A��|{��[-��kT�chx�"kUƑ�Rd݋J�xz~$LM�8a�����o���p)��:�@��������W�x�����pҳ�%���i�w#�Y����T��˯��Ղ=���v�U��E�օM��Iϝ7?��u}:��e;����?�^���������\$d��ԉ��#�x�q�Aq�����¢��y�>z$w����}��[KV*EXyzZ1rxƍ���Ѕ3������rJGeQSEK�
x��d�ј�t��",��jD@#0�,BP]�Ԏ+�{�o6B��`�# �Q	�b)��S?�S���"WC!a�� Q��&���?ޘ�����X|�g̃2�k!��5���� ���>q� "`%�2c�\�ϱ��|��5A#d�p���)��Y��SS��+�eq�1�Tx:�JMv7/��%��En��o��1x�z�|�9I!�90g>#8�g�{|�S��g\����B���9e�Ⱥ��`<��G!YۋX=S�G���Z�زѱX���oY�V��`q#�wQ�ԝa���>��v������*������/��/�JC�!�x�x��`կ�fk¦�&���.yOP���<�^��o���*a��\����zљX���^����?4<�س;�s��:d�`={�CC1`Y���Z)z��MDe=��c�n8�?�s?�.?��B���~��XlJӫs:�?��n����O�KZ�d����U31y���3J�
�T%��$��9"�����H&����c(e���0 ���AEW|Ndp|����P 
�i��5`�r<��#�M-�2��=W�.�����w�����( )60J���#^�Uv�@H�(M�8�l�(�h="�Sȱz�S�[�4z�tXk�����=I�r/�)�9�p�0#J� �o��o��������yQ<�Ng��k����_��1GY�o{����\?�Hyf��{�r�5xq�K0���<	�`�s���y�y�]�(1=9�$
��cC�A@�O�G�@Φ�A9�xm@ ����܌�{NOO���
+Vm��q�dDF1#O�n+#v�gdU�&����1o���|��Wݐ�6�}�q�;d{v�
��B��jՠ���(�:k����{����r�3=^�^�:�}�b8Od����zc�1�]8��kqC� ��ix�O'X+v<ȄU_�2UySS'�����0p<��(����TH� p�����1�(-.�⧥�5�_D@O���ܢ'C���R�Y<cˣjV�> �P�i��;q���o橬���4�F�^}��2E8���%�l�3���6m�����íJQ-fq��`�����)}!��CmJa����b��+���ڎg�}q�W��ann&ǳ!��ξ[�J�;,L�x����q�V$�	]�=�ɿ�ï���9��������y�A���=�;�U�R�+k5-��9���y"��b�f�i�0w<�>���|�Z��
k��Z�
n�[����0��۰�yF#c'�@��ŋ뱩{��J 7�2���pY���`y _w�e����ed)u��g4X��@�4O�si��SB��g��r���}7<����~-v��n��
�X�[���!k7c~8<�Q`�S6��i�k�"��[��X�0KY�(�#p:0oa����h�BL@D��|���\�N��"���`���	�F��h6�R��4��[:��7�*V��)+9�#��kVPQx����̊"A
D�CA��V�Q�@�nZѫ�p\�V�'������[]��-*�Z̬�
`���ôЌ����֐�"�b)l^�󋋲Ty�Z~�P�������R�(�9?����MF��5�y��&���-�����P�����Z�x)�/J઒5-@C��$kIy���=�	����ow8�,1�jyF2���b(Z��w�M�ܵ���}�㠪�j�Ra��,8�?���G�v�X��Gl��N��iv3�:ˈ��N砤����l6x.@�p�?Yh��T��5�����+�jPp혵�=�v�Ѻ��1�Í��P��r�Ki�)�G/��y��!��y���d����A���j<�bL�D�V��)
5���c�P�	$�xpP
��	:;�!qq	b��>��M�⽲p�������c;�՜
�aN���i`�x;�zv���]xͲ&�=�(�S��`u;'��~	�Џ,e�H��yT ���:�\|5�Q��
�Dɠ@eJ��V�J���_/�%��*���)%�YB[��g�yu:?�PE����=�L�e��6���C�{!������ҌyaĚ�b�I����Q�T=�Y�7��ҕE�̓��	?��c����x�<��=R��A��ʘ�:ԁ}����K���"����}V��<�F�!�9� ��e��8Vu����X��O���m�v�� �n��w�\�Gcü���±�v���/5�W}�x��5���� ���(v+�2��ky�������v�8����������)���[zo�¿'m�,@��b��kæ>f�\|�ՃU276aa�jU�
�j��D����h�pW5��R�X,l򾱪�_���zVi�X��nq��M!���`��)=�}��F9�@m�f&OXi .��/D��Sh��螮�E��@#���|QG�k�*S�*�,��զ�q*�9����ɛ,e��m��;�D������"v���)��M+��{A*���'˞���NQ�oR����b���GE��x_�E�:X/BP�|GN�R'SG�S�'�R�j1NDy��!6J֯��xMp�FZI���EV����hR7�Eʇ���}5�)��ސ��Q
�7<%��p]��ĝ�_ۧ[���Y��X��	����7u��k)V���O>Go\�)�궜W+�Y���;_~��Q�"xU2��A�P��z����X�p�I�8yȦf��h<{otl�O�ѵ�[���=��9���h ���@����R���/��pn�G�n���%��+�28d;.}��~t��{�q�/�ff	tl,l�Ma��p�[�v�?��Nz[F���f�0�ʀß�?15i>������ٙ\�a�PQ.4��m"��o|�]WT�2�,�Y�p.Ulr�aA&��ȐMM#`��מ�b�i�}1�SV�E�()V'㪱{,,Zܩ[.8F�E��+�@l��(�=J3��L��������"}F�KiR�Bp�vJ��ІO��H	�t^��8H�C
�A�Y-R0e����|�@�E��\1�w�	
c�W�R���~��`������`�y���2�39硃G쑇w�.���*e{�?~�cSk���H�կD�Gw���"{��̯����mϣ��z���|�n?)��������>�1���
�5V������e�:�������O�/,:�w@>��OL7��)�mv�m��T-�{�1��I;r��a����t�^�5��K-���$7zPTp���C�R经��e�����=�����<[�9���m�}K_�re��d�uY�-7�Ɩ�&���m������&�����1[j�K9��˟�\$C�v�؃>ܫ�A��-��ԜW��߻/X���۾u�W���;qrʭ%pU Ua]���X�XTy�)���"J3:XLT�����qZi�܂�:2��`�dn}7X1mk461�p� ()�V\�7����J����к�BM��x�J�����R:x���/O3�FA��6+E(+���N{3��oY��W^�g_��)�df���*�:��C�Ǩb7e�1��
 ާr�c��CV��`-f<[ɕg�6�
�Յ���k��u?~�F�3�{ ���Η���V��}�/�ۺ�B�Fl��v�ȉȔ�U�
B\�v���b�����dT�Ѷz�ӥ�LƐ|����>�����F�e��I����^���UNi;kW<�Z_fG�ǵ�v���~�F���9�m�sX4XV�?�a����A��X_4W%��q�I{##hn&�2�����߽�A�������
��@���:	�em,�����^�:aِ���??��C^��7�´]tA��k�� �`�S�@l	�
�C��7��qA���H���(�B�ě���<(�{��R��|d8(� ؏��a���SRb>Jc�����?��n��\8�(�J�U,E����<�y�.���LA�³�÷�>���r*���&�0��۶^l/���Ju�9���q!��Zf#m�?�On�(���`�K�*V��T����v�R�g|��mlt�6l����똚8�{��ͷ\���ꫮ���"�C�'���͹3b�\j��¿k}�8*�&����{��?������k~��ʾ�m��w\7`��G����#I�t�����
���l��A,86A$gY,-|DiZ.k�J��yN�<<6��I���U���������d=kA	�J��XP�Ƿn��XZ�J��uKД�F ��k��De�G, /��18<�4&R��_�k��)�f1l��L 7͒b�Aq�7���]r��8��ķ����e�(��Q�U��K�}%�Pu 1!Ȩ�`�/:<K/��m[!^�f$�9d�ʒ�1��_���;�3]��& �Eߨ��}�?�Ǐ����g��Ipu)��`OWka�+3G�nt��k��=����l�5�7��-+�ݬ{.�<>OL��ۯ�{������Ïtء����=g;y������I�G�9�!;v�����ĭ(.鞠/��%C�u�����ұJ6��4��[�5�UF*x+/X�,�i��a(ȉ%��R
�-����*2�_�5kW�f&X)��
��9�aSԃ��n�*�����Tc7�蚗=��������4&� �A�PP��5(jkՙ`m�D��&댵�\�X�.��F��J�e}��N�=�¿�c���0K$�TZ#�t�K�{Zl��S\p^uv����d�n5�Q�r�@��g�'K�Y�1̼�pMk���.��r�`���Vm�ӵe�c����50�}�@'=/�����S��?�u.1>��G��j��P�4sQ��I��f� >���ڱ#��Ѓ��[c��68�6"�Yg������{����X���=����Y/��^��0{��ĉS���7�Nǃٺu�kjR�H�"O��*�͡^���ȌtNh�y��M#r~�|Xboy�[���H�� �U��1���
k��M�)<�x|��a�u��bFbN I��,�X�|~|���.@�X���0������ e@!$ș'��
�2߅v +{.��9>� ���M9\T_����W�@V�����C���J�5-�c@l((�c�߷϶���^�ĩ���^��AI�'�
H12*��^ĐY�V�����=�����͆�K�[τx=x�����F�!�c�p�����s��/X�6OTP]C��J�#����z��:�@���l٘�L����p�=�e���C�r�������l'�~E^1x��ȐkV�W�?��a�~���9�m�k9g?��MF&@ڶN�����]'+@�N,!�m���)�,k��+ћ8�ųe�6�eu(��G���7i����N�5�_*���`�Ȳmx����J/L�۰�y~�|e�Ɉm�u�Ќ�M��^N��6��5mө5�{� A^�q�7�<^���C�����\����<&�@��7�f� ��@)��0g�S�
���O�U��b���=�sq�*�3{�{1���"ݼ���k�>lr[��0s�T����g�Ůt1[�*�B�p�{�3���&v"��稩�~p���磔g�~�����>�E�r0�����h�2yj��aϊ|p`8��`?�8<��
�sS���Mr�dYɺa�@[1�փ���j���E�r�������1��Qx��%� iǔ�*��HpG�l��6���w�c{}�S0�cp�K�c;�J&L:9���4����k��a��!V�z�:�8���EN�ų�b��HM��5�����Kҁ��-9�T���lԱ����w��e�h�^_�җz���80�x�"���5��]�g
Ͳ�T�+Д���u�*�4�3����C���H�lWk��y�[�nS��P��b�K��xz�Vu��<n���*�p��u���T:��xN�� �r�ʼ�T���^�y�{�{�.�(��^�w�N�)^)|�Yz ���P'��[���%#�F�sb&-�/fe�N�fy�_�b(o�EΆ�J�5p~�a��}U*8'�PV���uc.|�+5��+�A[�b�M�<n3��
�����T��F����ٯ���K�D8 �`�KR����T ȿE�&����`����վ��3��,��CL@5(	������{�;�5���u�`�°��\`�:7�Tf�F��\�I�~+�o��H��b�9{�A�_�i��[���!�2�T�����#�S/GM
�R�c���m�2h'��AM�u�����}�7�tP��*�3��ꭺ����n�"M&sJɤ���(�L�������}V�>ޅ��� o��B�4�Rʷ��B�"��&�%�M��w�����:�H���q&&��Z
Mͳ�x���݂c��^��ѷ3�g�V�^^�Ƿr�/Y���
_�W�g��r��_�,�aQD �U�+�Y���`}i
�x�u���f�ȏ��.<Y2�87q+���y>G�&s��L�}Z����������x-�̤>~�K�8���ڧ��e���]�:Ԥ�R(+A��	�P
���v�N�H!�L��lN�c�O��{:7= D�!�������E�O���7��_8�D����WK6O��0����yZ}��7��]b8S��X@,l�XNlB�(cH�/�>�g�8�ڝ�X���d��˙k�ͨ4��Ջ�Ƿ|�x1��@(L��Z-�9.�X΂!����W��pf	
�S,��ǎ�m����>���ń��k�����W�5}z�}�Mp��H��~��6^A ��@U��b�]�X��&p>C!��Q'/)��A,�Ua�|�T�(/��N%bX7p;�X��r�t��WD*Z�V��ͨ�ݓ�#6T�g�gڍ�^,+R�g�z��ݷ�H���߽UZּ%�P����t�z�_xB����|"i�����v��t*	_̕�,
����S�8��#v�P,D#�'6���I2O<�y
�,��<��m=�U#��ֿX31��h� B@�����x"|�|��e�� %��Y�+_��(��k�@���Y�{<a��+6!��6�|��VsQ@$�b�s.���!
׈��us}�n�����Ҍs��-K;3��GOZ������И՛���NKy�q_f��ќ��p$U���PBJWr�C��!�o��}��3K|���z�U\Z����Xe����HcbStr��f@���g����]�}�6[�SCT�5��>u�U1����6�)n�~�Db=G�f����0����!�	��u�]��?��?��yV[f��8�)�|:r���g�������:��Fŋ�,9��S`]#�	�-N@��MQbc哵�<$������ �`�������z!c;B�Nk{���hp�?�����;.��1}����=�R�
̺1�윘f��+���b�ǐ�#��Wa1͢��su��q?g����ȫi{č�ajh�*�Gd`��Pڨ�r^�q�[/\3X�O�ɩ��lLY�B5�y&C'�T�f�K����dXv���v�����������3��e�,TQ!���:R� �bS*R���pLΑz��-b7Q���[�kJ{�w�J��G����`G��Ҥŭ��BOEe =~�u��.�0�V'B�@si6;�6u����e60X�L��R����S��~�=��RA�������k�57bY�w�l�'����	�?װ���,��h����قֆ]�*%��!KFCʡ�i�����ڀ9�s�C�Ϯ/^���<�Y]7?f�0�Ώo�L	Q`���N����4ax|�C#ܜ����E�	^��#G���NT��GP7�L9.1+�C1CF|_�\���W���wߝ[�@TdqM�3S9�������A�F�+H=Uj��STM�E��t%��Ub_��`FE^�j^��ʱ~Wῢ_o�K������HcnE'Xd.�ã63W咳��ߙ�H�j��ɫ����N>�؇� Lɍ�?U��-��ۨp��[��0SL^V:̅w��OG��H����O�)O�,����}Ѻk�x� �
�B���Y�D�um�`�5\Ѵ��ULS��� �v���S��Vp$�oz�0���9�$2|=�,�_���9�r*X�_�S����y��A>�&�K �}@�Z�~�&c���d��yۮGq�PO`�� HU%��'q��a���"�H��b��z� �S:���ؗ�={zF2rZ�R?|���޵?Ҡt#����%��2`'NM؇>�1�[+q�r)ҳ��xj70�HNq���8�����kg2�S�]�W�-�ʧOg�*F�`۳^�zV���ز����L�X���l�b�\�X��Y�~]�y&n��CG\H�2m�~�r�����Gg��I�+���f+V(f����>� �o�^8ǅ��Ӷ�SǬ7PX0��N=��<}�X-x�j^㪻���ȩr{�4�$��M�et]�0�|��G�A������w<'�Y��H���� 8��n�B�N˶|�����/��҃8�T��� hUg�⫵���	��ˮ
U�9E^E���[n����҅#��������Kw,踆��ګ���^��<�)pn?CŇ��87^FJO�2>�q�t#́��S�/�#|�68j�����ÐPQ��������V'�g�M��Zu`>�P�j+8w��}�R/8�\��G%�u�!���2��G<@�j�1[Y<�kE)׃bf���E6��l�+J��7��g��/�������lm�-8�7�!�O��v�~}�T(	��8(���]Ps��AҎR�"�Ry�ί�"�Bvn��e���v�ѱ����63q�]ڊpڠ�����v��1�7Z��o!.��OC�~��2t}*����L�I$����jCҴ]�wޙ	^X��)e�T�3p����%Av��AoX���sX�@5�a�"`��w�ݟ�����?T��^���G��H��X�R��<� U ��Dv��Ӵh-�����xq����+����Z9�^.e��ю�9/�(��p��XYO��� F�������U�G��������>+���Ӿ@�(�;�V���W\��Ä�����{<��޻��yH�����Ԟ��:��'�Q�S�*�p�c��\�dd�^������	њ��K����6�zԖ���۷�'?���O�J�E�+���,���jv&�h�������~�� F��ќsvy�x���#v|�DX(4np��J����-"aQ�pN8��eC�Ñ�/���,n�w~<�!.~�������� G=��D�),�!/(��5��Y���<DV���])"Y�b��wxM���f��*૶�i���֑��hX�Bܣ[�;y�n-�:�Pj�~�]s�e��m�;
�v���ܲek�˷#)�"B1#���6��R��ѭr�s��
��`+3Ii���]��ee�n��Y�������;^���	�j4Ȣ[�n�]{�u��ؾ��/�}��i���a�I���^�{D��۞�^�^Y\���ӮZ�?3;ִ=t؎�<�^��Uk���>P# �����0H��{���ܕ�7X��>��O{���:�&���`��Z��ێa,��R��������U�"�x'+Z���w� �W��I.�b"K-��z�<e�S���^N�x^��d�H����~��7k�կ~�c�<?�J��@a�b�s^�5�)PSz֥:�!�H�T�#�X ����Z���Utυ,.E@�F���9׀' ,�aD��9�3V��?�)�Mk�i�,CZ�Qw�(f����Ms���l�����٘v��z��s��@�o�{,��(OJ��w-S������x�N瀋��	o�>�Т�
^��V�U\�ƾ��_��_��m0����U�7sYr���z����.��U�9v�O�S'�z���������}�P 2<4jW^y��t�-62�<�Ղ=�Y��Ŋ++���@Ѝ�����@�
�Op�~}���h�z�С����o�ӥz�A�"��l�s��^���^@7���\�;��3�"DbKq?��lY{jB�TF��.E����xr��M��`�eRk{��g�D	M��q8���{�oe舁�2(�3����Ӆ;B
c��Y�<w�8�a�C���j_P�b�NF� �C���"@�F
�O<asF��c��I����7�r�l�!Q�_��p��o���N���Vl��Q+6P�ᆗU�
h��Uʶ�.{�*k�>�2��̝���E����a�L��=�;�p�a�^{������g�|����m;l����-ۂ2\m������c�֌�ٛg����Ӈ��z�_����ş?��˯�ʞq�Mv��^���G�O���/�q�gT�6�d'�����^��9��%�@)da��*'X�����������{(ɮ�\x�[�s����F3#�r@�H��g�c��f9��᷍��l�1^^��<�m9'EF9k�&O��t��|���s�ۧk���i�3u��=]U7�{Ύ��6�<����je���Mo���IY�Rs�̝�d͊3L�U��et�������?�	xu1Sis Kt����o���`�ca�} 3ȹBW�
�=?�%�aB_�(���H�Q�.J���C"B�j@��ר0� A�
���8����y��F
! ��~���8g2?���*��_+}q]8<R�EeP0`�1��4X�^�O�Z ��������Bޜ\���n��f�sޠB�O-�N#tC���4��L�RN8�@�2U7b8�f!N8-�\G�n�e���O�s�(;�C�w0�Z{ը&O=��<��C�k�.��^�z@
ټK#r�����]���x�,Y�'���Q�������cn<Щ/��z�����JcґO�����X���e|b�P4�5K�Y�bqT���?��O��x���C��&�Nc��R��8L��$�Fֱk��X��C�����=%�܀���C��<��~�;9�6�ɪ%G�`4�^,�-@lѕ�H�
g
v'�5���k������=7�	�P1���;`�d!a���I��*]��� ���� � X��
�TL��H����9�]<�&X�P$x���964�EL����E�Dx��H 7���Nd,�b�sa����f��`դ�W�y�j�G����Xo{:�^'}�+͍���l\�Z�5V����`�5,6�D5�>�A�HO�ׅ(����6��R�A��1��wE��j�T+#�����HWg�Tj�תқM�T�.G����?�o򋷾NV�� �V�4E�o߷�Y�/£�4������4�X2`M���әH|�ټI'z�2ٻ���.�0g� d�'&�TQDr�h�/49�%,X���〛qO,v4u�{���bs���l� �U�������\WW��s]R�M��A�KJ�c�D8�U�E
n��K�5
8�t� ���%*��%� �c��AE�nPldN`C7��P�q~���a�@���j@b�x6pg��W<8'�)�>1�sM�"�����H$*$|��̑����)�	�m�b�i�G^S��Ϫ�*�CU��Ra�,{x��}Kep`��������S*X��Bz#n����Z+Y̽\.�1\�=z�GO ����U��ɸn|�P�z�>���^�v�^GE&ը�zGw��G��d�X�cE�_��l���39s�F��{���q-�)/�-�6��BQ+�V�IOW�.��F��$��QT+n�Z����,��`��,-kzՄ!����P:q�:��Z�܍ՔH����w�i�6�&Zp�4'�[J�$"��jm*!��u����ez�hm�|,a��.X��Wb����,m5�^ ������sI�8�/x��$�&�V3>%�����B4�����}�vZ�Q�!��i���W,�����J�|�FXc^ ����������a(�C�^=6��v|� �C�^j��](��ߧ7�VZ��Ĥ|�d�����T��	|��޺�e+�������·�#�x1w0���IÍgxp�n��s�:�3���ۗx�&9
������y�]�s���M�����c�V�ϼ��Z�S_��3�< &���C����
�:�L6�`�@b�V�,Zj�<>�)��vx����}���l������©N[s��UX�P�\-
�x�FT�D0
x:���E��~*0�7��ix�e��!Y,~��7(YI�CқL�m�ϳ;��v p��b!+�ɷ��h,�:E��!Zm��S��}�����>R�gx\��a ���&�}( �����8��7�zQ��(�ώv��U%1X��~�a{���G 
��f�}	�j��`�խ�5�=��-�S�խiz�܂��
����rV��� k^@���?�cy�[�j�-6�G.�=(?��֮6��e8�
:�!
J.�1T!
��+�*Γ���Ge��{�
��x)����@��#)W���V���|.)�w�>��^�x`���QmG��.'����Q�X9ࡀ��ݿ�8���˧��8>��J"[�#��ȡ]r����EK��j��Er
��"RQ��"�T�z��p�� ��A����	D�A��ˎ�c���T���2�7x>��b<|�B����]�Uxn�,~"�$�'����r�}?Nx����Yx�n�v�f  �K����
}	��N!\#'z�8P>���:������nB����?C��D�W*��K��uOEe��2���C��t�%|����6�~$�VUϿZ	�=��S��;�}�{���pohbO����"e�'=8���f;���T���CϛM �$��>�1'�*�(F�FOθ�f1���9�S^��4s��ɴn�j��X��8��o&r\aUh��x�u]p��@�,����x��K�\p@䰘QJ�67-Y=����=\5i�8�o�^ߤdԺ��"g��8H�X}GӖ�v�K`���0g1�5v\�\�>�*?XC��;=dȇ������=IZ�P\|nx�a�@��eX��C�/��&(4d�� � ���%+������u�p�����Q�Qt�B�v֔�|w�}��
��q���ճ���o��8��)����Uu	t�E"jm�z_wv�˹[/�J��*�T���O��_�.)���@٤Ru?���½c�c[%naZ~���?�01o].�V��~	5��ať*R*oV�[#Se��Z/����i��~�m�w�AV7+~���~�*[�H���'�L�w�v�Ly)tvYy�Χ��2v��i�+҈��G������w�y���w��][����f� !� �a��tv�?2�o�BKf�4�Ua��EO��?��B\x8����Z����`����2QeT�~�C>�>�n��,ߘr�J�g���b�����Ig@4
�:�g�BKPX�;P�q����hL��a�T�����60M�F�9i�wS��EE �z&e�8�9���U'`1���H�m=2�����,�G  ȥ ��#���!�t�2Y�j��Ke5�ft�ܪ��7�vmM���5�\��A�H��}�z !^.��������X��v���-MUd��{e�sd|�\x����'d|�l�7����V������(H\��7�� ����E ��<������q`M����z�굌��ş�2z��1�4T�hp]�J.Hjűw�q�.o6\u�<|�zX�،p����I\��'6:��yv����ρ
�O��sD��B���0D����������v[�x�X,#�^*��|����W��(8*&�휺�p����w��@���>�)�V(BDØ�g�ٱږl��
���˩�V��=�#vC�����C���0%z(#B��q���l+a��6{`I�Ž!���G>��%�5p�}�c�R��m�](���P�ꀾ� �Ī�e�Y��[&�;�-�$j	�=���
��?�8����s���A6�K�bz?�C���iY�f����*��2tx���&&F�d,�.Hhn�z��u��$<?b�L�b��� ��͞������&]w, +��?�����~N]��y�.�$��8Ir��K�\i�yZCjX�ӷ1/�5�����p�c�(6g5j;����$.��a�ǯ�3���%a>O˟�B�,c�8�6"餱|��iE`�g
��(?���{���!A���Y?�����-�F/�`���U}�X=�%r�Tn�}p�O�Tq����L�#\w�QC�� �_��_J��0ҡ�$l֧� 4��u���Kj��a��AȝBΘ�׆36�5��h�ò����C�䓻��-���Fr�q���uq��>�e3/�FY��? _����u��U�rM]���iG<p׮r��ak�GͰ^��Ns)�q�C��p<��|�3�7�Ɋd �#�V�+^�
��W�l^+�i]�ӗO�v|R'��dCv=�CjU��֝��@>+�5���E-�T:�����Xp+�%��'(F�W�p�P���'��yQ��µ6����0"�Ճ9gXe����e2lCd�X��7C/[�Z�:��q|&*B;1��҇g�d-�E ���Bx#�okk�81i��By��l��R@�*Ž�F�#m\�į �݃Ec#�q���ڄd<�1�E:e׳~
4϶XQ��������A��0�BD(��Ї>��ϸ�gp�DZ]�{�!�6�����J]��d��@�����<8j�����l�v�z,��� %�m�}�d��5�i(x�q��V#p�bb�(����N)td�%/y��k9Ier�eW�Y��&IN6��*�U�����1w�?�c8tP����ֹ���k���H�R�����k������X��Q���]ۤ�_j�Ѓw�#�X*�:�gƅ��J@%�d�.�?�.�@�a�<����r���ܡ��pNl �5躓��վ�L����7��S����?���~׬Z]S�@y& Q�=6z̅�j�%䦳7ʅl3c�;`�j(�񊅐�� &�>rԎ�Y�0�rd�����{l=�
7(�8��EBki��a����V����P 𤡸 ��}�8�����Xƫ�Є�f��ի��[��FR>�����è��F�[^�R�3%5�r�K�������ռ�`<��/���y9�c�~�<����84��+��I.[-����\�(�~��!�c`rtJ>����C�<x\�x�(l���s�J���}�0�x0�L���p��T&�~��񉒹��t`�@�����pb�@� ɋ��x<,�~c��*!��.#,�|v&_���6���ŴI7hd! @��
S
�C���,,*�zc���D�c���  �ň\Y+`�!,�{D����m�/n�ه�an���<��>{H�;M�	�i�3��:,rҋ�w�e��_�m�ug�  q���7|���Hр�`]�<�'�>�{"�k�9(!��\ӣ���v`|8+W,�m�oAה��!�`�aF&U�wu�[���j7xwu0���$���ɸ�g쇛~��O~��	����J���M@�Q �	��,�[�J���$U,tv�cO<n��@A��!_0׋Aӝ��?��e؇}E��"��K�я~Ԅ?�
؜�dY��H� Ə���b3zǬ>,�?��?�ςW�f�|�4��bq�����gB��⛵:�B�T�'Tk	-��h�`Ψ�Q��m��CH���j���.�s/ ,0Z��� H�`�ạ�|b7Ɗ�����i|ZgZ�0&��� 7���7�O饢0	��[�����ǏkA��A��w�wm���_��	i6H��>��4��:X5�A�c���뿶�!��ϡ�PQ;T���&[�c���9���i�5b�sd^���p*�^�Z������\���s��z�"�^�|Y�|�]���S���j�Q����|����8��q����D����d��/����b��)/��d#$d.2�Ҙ`,>L>�U0�c��7,J��ȊȒo�ƳM#�}>�O��C�~��`�����;?��D]E��=$��b�r�@#�nD�"����C��Q5��mm9���h%B�����_h����{��d
d��j���XD^��/��`g)���>�|����h���a�\ ��{�]���a,����`������8'�C�<�������ll�C>�=7�R�,�FՅ�@��ϲ�{�T�޾���⹌�=��F	��� �R�*ܔz���?���9E�0����������=<G(W��^ �'�7�1�02�9������:��|�5~r��˰i�4�7��eec���Y���������0��I��k0�E�&�	�釞����EuH�<��s��0���Ca�L���U��2��m�ԋ��&|��ZG�o������m����Hos�~��o�+��aeb�A�����p,��/�.,�w��]	���!�������c���#$�Bˇz�ӦWɦG����i���<����M���Y=�U�@���7��ֿg���۴Y���K��[R���*�S���64�JK-UK���~��Y�HH�sG�������C���O����-���bIVi3�@�EzrW ��S^��7�Z�/Fg��������d�9��O���,6,�>�$P��d �Gr�%����o��L��:J�;��뒎�ZS�qݼ�p�k�}#���:�7��!��	��[�J ���Φ����>.��8�AC�\�X#C2n����7���a"EaϺV���%��3Ɍc5�c��B�'`�1@t�F�*����A�ǳR����'���w�Q��f?3�Dm�r��V�4�����m�:�+ӎ�>�0}d���������w[��Ph��½HXã�L���C��DC
���3f(��c���c��b�i/�1�L\{̰�9>���
�Ho��\�x�X�
��P ���U���[� V5?ϟ�l��l}���oTC)N�%�B��KnNʕI��fBG�4R�ؑ�ſӨ��F����n��D-�b!j��LaDWߧh�����rV���X}�(r�P �*��q\*,����J���P��	M�@������@1�G\��J��%��ҟ�]7Ce� <�??�R肇�ew��fA��y�汦,\j�9�_��P��q��=�1�"(?�opݸ�}�c���7�5��"�3�O���lY$��>�~=A+l�?N_��<��R�\Z�\d~۷Z���9c�<-��H�!��W.x,j|�)3�˦|�87,�Z�YS�	� ��e�?��q�wa'�L�l���j(�0� �AT!�,F�i9?l��>e,�n?&;�:k��(��!�?��}( h�0�DCk�	��6\��!b�T4P��nR�!1��3�l��ռG�Q��8��CD>�r����Hv�V���!��c�L�d��P8a���֫�7���q�?�9~��=����?��$J���L`ؓρ�<�$������<��fΆ������Nߘ�|�_�>'6�o��	�kCDxDJPX�'j  �a ���[@̵i�$�oq̮�&�՛����~�)�nE
9wO�c��6E��[D���,��FvōG+�����s��%�[t�3n���R{,l�����/���6��/0(�0����g���}�LBC�x��|H?��?�Z�~�����ѐ	F�/s]��ܵ.\�а��Z��n�\V�"0@�{F�����2�t�q�)��2K��h�^)ǐ�ؓͪ�E�\<Yw]4����	��g��)�i(����7&������':N{����;���VN�oՐۃ
�V�����	��l��e�p� I?"�=�S��Q� ��PO���ftb�^�D�T���F����9c���;�q2G�e��o�QPxFC̅w�1��\���;(MT�T��F���#�?$�HoϠ�^�A�U5�O(N��%��f��	z�T�����"bh�ъ��|N�"�@Z�E���IfB&9�,�ހ��i��!Z/P���s����T*�w�voeA7����r��n]��DTܗ���V��Cf�l����� �Q7��@7�Q6��+Z~�M{<W��kQ-q���ټL�F����K��ua�Fv���9cI^�74tHB$��h�3�O�"�3iT��4ʡ�-�8��a蘈?�C3ĕ��Ӝ�8��|��ӧn�`�#Q+��LK����f��|r�3yǇ��{<�}����ύ�$�,����T&[z�r�H9��(t��
c��b@Ӏ|�]}�cm��8�cv#��]����n���o88rW�Z:���V�e]]0ҜYŔ�4 %p�l���}�*x��"F߈�	^�b�:��̣�8i���"=�٨���4����  ޘ-.��Td8�w�h��°-v��|<.CA�|~a?��\�KK�_�R�ԪGb\+Y �b��Ѐ�Ti��LUʒ�,>ZE�_��u� �'���Ӷ���6f�I��v�t���)[S&4a�u>U�X�s���|Q[H��ܴ�vh��˷�����'8� �a�Ic�0�I �oȠtj�{��TP �L�_?Q�[��<O'2Ny�?''r<U���3���	.�����Xt�(�}aތv���Wr0���#�J�xD��k�f\%��
�TC,�+99U�kba������7Bc\�f��Ԙl&������h��5Z�HrhX�rprj�5H䆇G��Iވ���d�*Z.�^�W\_$v��'KR����d&�l͠��p�&�g�f�0����~Q��_X���F���?�8��f��%N�D
pChd�3�A�؊�������a�M<N
O�]��Dt��&u����bh)���D[��{��T,�F(�uߨ98_�~�]����I4��26Q�#G'��k��ϿVV�X�\/��M��'{�Ʊ1�T��w:�����ό�J��zcK]��K�O�I�Z3�P+�Z�
��:T�ҥY�'P�����U2Ĝ+:K��x���]�`}�^����V�Npq�fU��F�m˿����� T��1�6�\�p��er��73X��&�7M����y��կqpb��)Q�ҝcl��u�`Xv�6�Å!:ؔ��y����ʰD�8��1��;��T2k��U��C����%/�ŘH��5��7�~'�W�q<܁Mb���dE��>�d!�	��A�h��Ȯ��Lޗ��I1P�g�t�������6湟�;��u����毙�ol�56wMM�y�Ӵ���<���6&*����<�Y�ef/^����Le�4,z��Ҥ|���_��~/e��W�6?�/��[�o�Z1A福u?�@��1�f(�����8P��`�.�#�����d�gZ!�o�:����ϒ+.�\���oX%1��(�:����x�Є�iZ] ������U����'�z����1{9�r �=}�d`�Y��=�׼V�{�L	�(+��u�Ԫ�U���#�
�Ը�FG��L�wMi�Fdx��f#2%e���;W�V��b���d�X��K�����G��^3���
�f:���2��%�Gk@@4*��<���(x;���T��3�!�V�7{���ǧ�f3�ڨV�,�0��,��V�..�!"q>���n�.m>%g^Ohg�3FH�7�����$��$�%J�e�&��I��H�V^q򨤲*X¼Y��;0��E�S.H�����y�����y�E�P�J�)r�/Z���@��@?�D=Bz@�`/�3�Z�l\n&�c�PF?�FG9mI}�&�׆�J@�����u��<Fz��?�����"_E�������Ƌ��c J�JY3p��L��z,E��V�?,GF�4b��.3�4�'��(X����Z���L[��D������7��g2Xc�$��|�͇tC	ԬaRl��=i^X3���X�˰k!�]������(��aPV6tx�>�d�R��R��Ȧ�Ζ�k�[�� ��ߡ1�N�E��E^QԂ��r�
\;����*��ꄏZ��O���k�����I���/�X�ٲU��XeM���j�`e� �h�fO,�׽�u��YD���ˇM��D��d�"����0b�ȬE�o�,��}��45i:������czh>��kL�h�!�'%&TL(�@d�d:�_u�?2��@������4Bm���7��u��b�/�G7r���w�h/��y����HP��JkB�}&��#'\U���&�èG@��g2ܚm4 �.���\�}P3u`-��}���~?��*��ç�-���	BrhP
�j�|̏��X�7l��Q�h��dVn΄P�2���Ϫ������ร�_��-�E�Е+_M�=�x��GT���8~E�F�u0.�鄷	^���GS�h�X�O+Q*��8�c��T��p����}g�/���(�}�1t�1�U����T'z0'&N����ȇE�?�}��(䬝㱣#*�'�|\�������q�9r�ŗ��3j����?޾=!������u:7po阡�I� [��u�\�|��pJr�H���%w��=����K�汪�h�����^����L}@Xl7�|�qsӊ�5 �>r�B�;���<����_�z����[,c�� oj�+����Mق���"I�b¬h4��E����&������|�=��A��t#����ZY��U�(̙�`a3��1��V]qI�zL��n8P��YG��7h՗a�=4�?	��x�e���sq3�,��~���5,����F�	�Oڊ�,~��±��	Ⱖ�جi"OƦ/tmQ���҈��A6gE;
�nK����������R��G�� U�j���5m�tʅ$Cԩ��~=����P�t��$���g�W�<AJ�����v���,O^#�a���$�3��E�Y�<f��;N83��0%Qz����Y�C���k�5FS�����@oP���������߃�����7!{�<!�|ر�I+P��p�9,O��>����] ��Ke͚U�8��'w<������I�)/�[�}�[M��<O7�9��f�c�%���[�˭��"F8:<l�����_Z���{�g�a���2��6l��.���P�o����Qs�����o���a���d%8O���>� ��:�ıZ`Q�*�'�N�B�gI�,�����QF�$�Z��W��I��.����P�V���<��*��n�JY��B��9"ׂ̡�G+�!�{� �Z��j2�|H�S�:�[��j}DJ�q��(�5e���;oT��Vc�!��]X�8_Ը�(;u�"�%�!�jჷV�U��KO�R����E�*m��N��`mG�0�9*�ָ�U^�q�:�*@Gꗊ��Gus#�l�r΀���V%�����U3�d�ff
�|>Ãa��-�Vፐ_:t�j�ٺ9NVV��6���
��e�u��ީVc~��ǯWFr-�����Y��>��"��L�����`���"��_��������@��=����j܌���!��I]�����3��(�՛�*���-�7��笁;d���0W��
~�S^�����q�s&��͛�ڄ���ʷ��e�ֳ�uk����	�6fdl|B����	�y�u�]g� x�Gy$�h�F̎�V�h,�p��2f�����2�(�}S*�U�,D"�j�J�B4�=I�f�E+{���M��5 �j:���F�4�.<�r���g�/��Jy��+׮P!1�B<vC�p^�:@���ty�*���q����խ���C~�
��� E{��321Z6�epi���,Q-���+��v=.���p�K�8�B;+K���a�H��UUL��0p���T,)it˝j�g����#�^�#�s�'���/�;������REcޢ�wthJ���άtvAY�1<�I��g6�#E}��[��u�ͥ��)�� ϰ&��f&k��,��nTu9z����O�9<t����N��~,������cR���r>��I{,�1`U}cF�k_l����8b.�Ǽ�����n�[ �B���z�{�k�;�������=�\�T����񈮑��Y�D��)kh?Uv��K��������;�'+V���/���m�'���>�ih�e�<兿��� ���U�;�Q�������q:\(&�l-�p��B�S-�1k�v�-��%�Nm�����	�^ U��݋�/��/��@7%߭$wG3�ۉ�f:�f��E��I�m�ΕMg�։�������*�.�_7�V��@U��C�F�;������b�'��R#�.�ۈ�#uRy+V{��G��w���뮽J��ҮQ7�5��Z�D�#�������wn����u�Y�e�:U&�di����*��>V�o�^��(ʍ�]%}��t�۰�W#���kBqa�'Z&Ǝɒ%r��W�v^ ���\�>�HY�ꍤ��Bjt����#�ߴ������*.T���W���[=� �8�s5>V�o|�G��^p��?�i�/��!��IC�c�׳����m�,W^u���Y�9���	�F��R1���}Xʓr��[d��:?u����[�}ʱ��7��GF�^���K����<��E�����0���V��O2|�B�������~�+v.th����Д �������#r9C�航���xTe�r�?��q:R��2/}�K���蓣:Gw��r�%W�~h�ʕ�������f$���k1Ny�ߒ�'r�-Xh��Uj�8p�ڿ�P��֩��::T"n��*�qO
ZZ"����H%
��;�y�?��/ؿ	�d���\�6�
�|/c�O3���#maX)(�)�&�,*��zք�6>Si | lr����VQ��ch��k��"��Q�o���@Za������MB�%��e�S1���ʢ�	ز*�@/���`��-��p�f�︡�
�M)XE����q��B!{p���Y�5w��]C e@��oOA����Gz�s"��a�,C�j��u�A��~�
���B��Tծ6�BөF$��6�8!�Qu�"2�IxO�������Kh�fG��(���e3h2��zQY��	bNcsGx����p�0����@	�z���Hf��q��b�q3RH���kD������F$�eMJ6������L( �u���
�9��!t!C�^�7 �@����/����jҮbxl|D��R}�i[��a��	�$��󙔮�kk�DgGo���:�q����o;�����Y��h��8D���ߑ�!>��x8��@1��o�����P2l���|/����Ic4[K��ɒd�ŵk�yF9�؂��'"5WSV6m(���+"6mEh%�w ��<F�v�C@�@�{�X]��Z��[,��>+��Q$�1��	,$N+�)��ͨ�"1�#�آ�N@:�G�a��į��\�ؘ�rQ�6*��UХ$��}�*$�E*v�Z�b�]U,���M�EU�����nT$V 4K����ҁU7!�S��͍����`���K��T�~�
�|���ME�Y�Q�nM|`������*�lƞc��C��)�C�-}h�':ȕJS�iK�?_���3H�\�F�"�i�0��.Yh{*c���ײ�D�I�;K�B'��b�'
}�A`�{�{����ޒ��?��^�*���lﳾ�͎X=��Z2��^!��kA-i�$���&��,��`^\�:��n�2��3P�Tͪ&�R)���>�.�	F��	���v+�5	:eCnQb��+-g%=<�^z������7-.�������/}�K���`˾���}�9Z:���9�9Z)��,�kp/q�˨��E��*��:W�Ѕ�`� �Ě���3b��#��Аad �g"V["^\6��x,���5�Q�)�@b��0F��s�H��0��$���g�TW��6��nө72U���В�����d�D���x��A�ϪL��.�	(�sʚ�l?D筼���E�(��'	q�!Y=^�����2錛�c*劕j��	{�~Y�5m	_�S�u��z�����\C)�)���=8�qEP�_#w�$�[�<s-�~�O��a�Cj��:m�P�r�����Fw�>!�Hp߰�Br�gfM��c�Ν������oΫ����q���8�RdH�l��F�*U5�
�NWcr``�<f����=.'�E?����?�@U`GgA�����Kz�j���V�[�{���Y#���L��DE��V����6����^ ,�������K��+���|�#����\@$��U�ܠz�6}͌��۳5��������B�)uOIU���`�Y*X�CG�&�!���F"��F�j9v���\�g �[�`�a�NQ֡�fE̽��N����D�����>��g��ʆH*������g����1�u�������]����%a������5�Vv���W��UG��r�p��BcYU�cG�z�D/�`�����16Z���^��;t�����|%e-���hk�3��8����
Wmj�Gz�X��$�#g)�JU+�����̑#Cv{� B38�SQ������U��l~�z-׀�9S^z�\u�T&&;,��/��B������wK?��Sjh��W�hG�L�2#'��ǖ�+����q��gn=�Ċ�0�^��D w��;��p��� ��?k�~���uk7ȡ�g���V�����n���~����I)�|��[^���zpL'ͫX�8�$�%aN��54я�s�v��7�+�-W_�y��{���.��]�K,|�u�u�M[Wv�aX�F�W낯�ӟ����P7�t���o���0�~s�"7�$�o��o���E鉺-� p���b���˖���:Y�|�)��v>)�?-S��%E��EY+r��`�2Y�~��%�?�^FT��ԣ���c,�L�
�^������;e��5�v��1cC>�o�ZS%#��d:,�X�5 �*��'�fQ-[�Tϻ֊���{Z���%�)�\R9C� {_l7��8,��@��߰BV�Z/�� ���'ǆ����,T�kjD����������2A�D歹�T �-Y�v>*��~R�"ٲ%�%U�L>�)� B�%�ӻB֯9[ϻN��1����U>�T����K>�ڂ�)���\��Ⱥ���Ы����?�C�ј���p���R4�����}:��e�ʵ����d����Ԩ	�P�	sVL('t��Pa?�B�]+T���9����^��\6{MHDW��؈��4k�DӍ��j�}�8��1�.��ϱc�~��_��_���E�@����Rٹ�aٷ��Շt��V+��;��e��~y��'u�����,�F��@~ͼQim�EQx��}��#
m��bR�㮻�˥_&�j�#q�~�9rdhL���'�ʭ�1n�p�W˦�ےb�{��\>Ұ����`�����|�k_��Sf��1��s5��q�-�GN|D�C=!6�I�Z�Thde�곥�g�
�N�9��aCڬ��#G��sm�����L�����9c�f�����W�궚
c��Cf����X��D��2��@ϹV֮ۨ�YH�3Ղ�{߯
V��%��q�����w��sW��X-����JU��U9��rŹ�, ��^��N���M�.TA![P�Vz�d�؈^g�u���oZYU+W�wْ�r��3�"�ϓ�*��� @�*F��Qv�O*g�w����z7���*A���;/��R�Z������Wb�@1V��~�w�Z�)Y��G�?'?�~�
"�ʺ�v�zC׬�?��/���v�U��4 1ͫE�~c�����x<nq��-8�A� }Fh�۷\�:{�z =�,;{d�*���wD�1m��P�5Pn4�T��I����ǯ�hQ+Xf���]�z�z���~�����Χ���5�y�����}�3 ��[���!� $���սT���(���W	dr��Tv��~�U��s�7�h�Ȱ
�$\dJ��1:s�Q�Mҭ��#�������E/ԍ���^)W\q�Z~=�l���[�����.6K�/~�f���H�7��|�r�ԧ>eP:|�w~�w���a[��,�&�n!h.6���.���A�U�ꆯ��4fbq�n������.��YQV�ZŹ��~��4\��b��,��IIO�r�n�ֈɺ ��(O��c!�jC�Z�pܜ�TEܻ_��B-�^�2��M�b�UƻU��ˤ����T������Wk+��2���:u�;:���c&�sªY��l�*1�x����kM�@L��V]�� ����4mJ�����0�TC�W��֯�"#c���ڛD�4��F̀M���):O%��"�*�^�R\����H�`���z�=�dD�j�58�ӈg;Σ�s��J��Y��jYv�K�=�d�>��S%QO�1�U�T�w}E.o��z���Md�h�=�R�3�@�!��3:��~���X�L�
�Azy��y��F��Ac���%�F��<�P"�x��<�b�WR��q��Ss�2,tp}϶��ׂ�IՀC�����?���z��PBr�礝��<~Ȋ׼���[��,]��y���}�?�Ò����r�5�ɖsϓ��X���>�_�)����e�����?j%�<��U�� G�O"����)/��Fc�V���kn0aE�Sk'�ﰅ`t�z� �	d�X�@�� �9T��;��~�#y���-+W��!@iU,􁲦�O�2>Y_��X��<��,�zF^���e_'�ͤU�Bh�^��
��7�u����׾c������j��q�*���U2e�6�I�KRQ����m��yz�nٳg�\r�r����E��`�U`���{���&J�Id�����˱�1y�^��?_�EQ�mJ��
�@�W��MDQά�~���^��]�����ea�[o�U�٣Ϸd��(*������yq��n9g�6����S;���[/���&Y�r�Z��l��.[c��)��`�U��7�\6o�P��|�;ߖ��k����s6� �2B2��&�`EYl��h�֨�c�paC��?���ۥ�җ�D��id�t�B����*r5j��]{�z]c��#����9�\ 7��")輢�"�Ϲϫ�����R]��.ٲ�K�~�K_�b��oy�іXD�i��_��z��]��D�r	�^Bk�C?�ӞY��î}&@�R ,�\�
}�pѡ�:��S����ȵE��>X`����@fpO���� Q���A��k��P���s�̳Αo�9�������iN��d�$w�u��w�vɫq�~�1��g�o��=MNy�H+Ӡ�����y)����|�2Zg�;� �����N��z��g�����.��� ��g�/$w�	�C�ŀ�x�Ï>��lC�a,Z�-��8��%��	�@����Y#֟c��� �DW�j9��F������r>2<)˗ʹ[/�u�W� ,��ZX�g���Q��t�jA����19phH��v�
��,TS�ؽ
�2b��4�,H��D5�9����e�X��.�B�ظV��}��rV��87��0��eЩ2��Uo�wTWJ�l��X��b �ƘP:��0|Y��2}�y��'Գ�+�ܢ�|�����Vv=�A�!��"Jg����S�6WeAP6��@t��X�X(-g�EC(�]w�t� -�>�J����BY��K�QŠ�H2#4�0�Td��U�۷B��T{r���?d��\v��5�B���<G�0���e��Y�"/G����[^�U6��Y�*�.�Y�8�"��!��ݳD�Z�z+Crtx��vδyH�a�#w���q�.V�������9�p�ؓd�D�Ίeˍ��!_|�W0 �
�0��rYX���W\j�H��;�����s��##���ʑo盦T��;t�M�1WP˜^��K�<�pp������Mem~��ߕG}��;V�Yia��jo�;'���wВ�۷ߗ^r{�!0v��8>��Z%0*{�0�)|�S�4�Pr瓆�ս�	o��<���j���f�	*#n�r	N��']B�^u�!�9���㐁�$2N]-�RmqC�����@,�6�Ej�Ud�h+��JĪw+�X!mU�)K�A0cn�F;²�LNLY���c��ڋ�W����jgü�[��l�f��A�r��>���9���}��҃Ŗ
�"oČ��Ɋ	U��1cNZ�8�\6o���*5�r&x�:�]�H#�� �',i��@11��h��C�P!]��˲���c�5㺪��X>��Ƚ�T� }�g4:6ay�FX����n(��Q���x��F07C��y��F�,�B��R��ks�deGGg�9|�L~(R��=:iV�Ɛ�(YL������>"�"�P��8�~�Ϳjt ���� �9�����Y�c�+�
|�+_��M�e��.Dɶ�!Tv�ܽ��ͷ�q��ۿ�h��ET*1P�1�ZgA�����.�
���"&��V t��
�q��׿f�<�:� �U����x����ZR�0��i�� Uox������k֭�߻ݒ>��� �/��/m��B�G�����E<F��b�%����͊�@�WtE7i��8��u��L�"���$q²��nk�ё�!�mxR;G�GIP���0�՚��;��B](	�x�{n}"ǜ�U�?.	Cᙕ�QRp���¸f�Op^��
N��������g�{�.�7N�ȑU�K7�y+�r��(�M�TP�������I�0ra���Ūa]���)?\c*��Z��t�
�i�hV��P˭jJ7g�s�X�*�1Q��-����F��rE]��F��%��I$K5tךN�cZr��A �2����m�y_4��i����Z��>L�r?��e@=�?~ߟ�
X7d�>�Ʒ�������>A`㻀h�3�l��`�=�z]�o4��5BX00-�{�-	�#g\�l�m�>�[��X��c�R?RO,k��uu��B��[�(�B��׿�����`0"��'4>ڴ�9��2��2�4����a���&�1�npΨ� 4��̊h#$R��>.�g2nz��������n.X_��������/����!��^ ��@k�����2I�)�K$�`(���>��D">����2τ���["�P�g�OX��ݜ�*DQҎtnn)Zˁ	m�1 �,����"b6�~^㣅���ʙ�U�m��3�<S>������ߟ�� ���>�9�� ���D�^Ƴd�ܽ#�����T8'�|8h���s��6��aʹˎ!�3��Ȋ���ݴX	�B> E]�Ї�w����躄M'pY��\W���~�17]�t�O{ܪ�Y84�No|&:_���{Z��k��5$>����54�H�s��b�3���b�}2�{籉�'j�J���G�h���量>�-��AZp&�G�b�mmb�B�`O=�>��>�k����}�'��Z�v�F�욟04��W's�s�<�,��:�+rv�x ��>�,9�0|zOT4Xg8����|��8�k>�|�M��40��P���zh�aa�+`����O��L�=Sc�{&i-S�(Y��s�P8aP���rS(���>-5�"�{���M���~��;�w)l}�#T���y|AO��S���Ӓ'j������ p��2!Tدi~�|^�5�3�p[H�p<�ab��B��ÿ���.�G>������yoD�  b���-/ �
^��,����Ƃ� ��c����hNFs,�����ɤ7�'�m�i�yc�Vڇ?�a����}�����͍�>������7�s���P��L!�6�/�}�I���'��Mkʷ�\«��"6Z��5҂Ǳ���hnxc��y_�ӛ�s$�Wz$ �W����d(�a)���򇉀�����2���sH͖�o����}�~Z$H�4?,⯋VU긎�DyF~�g���-'k�f��u�w��N^��#��yDU?��y��ו�W�>���4p���q����O�
�h�%��Z9=c��
[�M<<�������>p�xA�#�e�^ ��6|Z�'{���!����+Z0��Z}��D�-�wz�x�gU�|�<���r��js�z|���|___b�3�G�L�B��p���A9Vw����������\�����4�3ŵ���yzE�Z����q�B�
�G����g���O:8�4p0'�(j��Q���ż�Y��+Þ�������9�=��Z�4<V��6�ۉ@�hٙ���Xsq/��/f��_d�6`% �	�I<
��M�\�}ف*e
!*1ߺa��0U4� �.9|d(&�j�X�͞�h���	�5�����c�3���5�y����=2|Ԅ�/����A�{�@b_���{�6L76�o��:g���Ő_�`}߁�"�s�u�b뉰�ߙ��@@�Ч���5%Z����>�(]�������-,��c226*ݽ=��:p�����87���8�x�~���:������>�~�]Ιڢ�c��:��,����Q"�S��[��g�dz���a��k��c��h�y��j��Kn$n�<^�uIRaa�c0AI4r���'�]��� �}�In��7�Ip�����l$b����L�����hY�@K���b��ap�O~�3�r4�f�Oa���.U�B��U���3ă�
!��.`�Y�CagB ���x0����܎�s��)�}t�����ߏ�7���00�Al߾݊S�5@1c#oT��n�5����2����s�d3��*w>_*zz����yP���<=��Ѝ�Ȍ��}���h�Od������ډ��L�Ml��+�u˗��Ń��H��p6)�
y�)q^�8�no��	&?]|�~8p�\�/?�����8�މz&�p�΃��_&�y���jm��9?��G��������ix��G�c���Ƿ���l(��0�
��6p�L��a���OC�
��Nǟ+*Z�;<��;���i�%Iq�A�`��V�)�4�4jq_+6#Qb�"�/�3hm>�� h�Rc��e�_�ͮ��<%]=�I�̚�x�]Za�d`�b�۱�ߌ~���Lt"j��h��76b�� 
����Ď,��~T*�d���;�8���<zܒMq��k1��s�a�#���?b��0����%T�I &�zg耉A?�K���R�;3|�����{)��x�����G��|�|��W�6س� �ņ�Oy�?Ο�/^̔_p�lݺU�����gYSr��!������S;-�%��'>���F�{��x��]���+
�V{��s{�'�g��3�G�{m !g�
D��oȽ�w�}VD�y�o���>Aˬ�ʳٔL��I�?/<���u����љ�Ze������p�g�s�>tD���;��"y���70�1�D�0��dCD����G{�������ʬ{1���g�^�k�J��_h�a�Zy���#i�a`":1��׹�|����i���J!!iֿ8��/|�M8NWwG�Ks! s����@ׯ_/o}�[�c��ii�~���Cdh��t�~���¥����h��h=f#h$z��믗[n���	�@0�g��-[�X��Aw�u�) �*,��Ny�ߘ��
`jr�������w�g�nk��{�N�x�K�ʦ�g�E�\f��(�B�6@�|�I+��
������_~����G�h_}�7�Bb�l��h��6RG4ú적~�K^�dFz{�L^ �������ADa��A��W��UV=��������F���
9�A����W_)��21>"#��r�]w�~U H����DL�<!�<|�zc�o��Tڈ�n��K����J�/}�|�ߴn^����jU�h�N���NȘ��o��h���O�3��W�C���GOW����ܿG����㏘G��R(�#����\x��&Pdx���lE��n�8b���Qs����s�\t�����)�V�etx�H�\����4���l-�j�>����ɫo�o���E\(w�q�'&�T���_ϻ�
��G��*��l;�<y�������޹K����h
 Z��H kBҎ��Vc���^'g�`�͓B}�g��^�23�ц!�B7t���o�Ċ��Rq�%�ʚU��V-�qZ�����cCOKg�*ݝ���RW����DE���w��񆛭��ٛ6�k�<��&�|���*�����o5l�!̢�}��_�ݲ՚z䳁<p�vY��G�ذR���ɤ�Z�i�6���P�~\?[S�������ꪫl1��G��6$�B^�}�{���7�2'�3���e�k��h�>�0靣;���Y�- r0������mo3��=��h�CV`�W+E��أ*+�j .�]�G%�	\߈L��O��ب�i����++V�1�Б����,>�:=Q�S^���a1�C���ի�J�^5�s�S�f������J��Svr������ݵk��t�M�;�Z��v[R��&ޯx�+l� ��\>(P=ca���( j��o��x��3�>��C�7�7I#R����W~�W����}��=],����<��òn�2�~���J:$�=-wv����49w�6k�y�g��e+�����/����-�g�
_8K��T0�)�I�VD[ɻ�O�oe�֤�!�0m�ᒱ*Z�����xa1@�Ӫ���+��������ϟ�V�!IZ{�G{���
\둃��;o������9~�������x����qR�<�{X����+�FJDVƋS�C�\iX��{�Tt�=?�W���Vk�T�K�Z��c!!�S^�A넯�42�M���{�|�;�J�h۵�C[?�'����/ ����/[|n����>=�y�<�$vj'|O�A�.l�9��G���>��gL��;�A�S�oذ��;�������-~~X�4�l�֟�0D���dJ��L8ցj��EǏ���	�5�Ԩ���,j�'lT+K��2����ٙ��֟4���0N�0H'�Ux��ĉ=8Y�����q�Xxn"�?2��]w��C�����0��h��;��Qx���ַ�%��ޝ���T�-oy�y�0����]�ش�'��P�̎�!'��Xod�4ʖOѤ�#�$�I�����r#�N�"�(j͞��4Y���ʥK,�a��R�Eƪ�J�%�q�1�ή��d�>�B�%~H�X����������\>򑏘�G�7�����Ѭ�����sj��>�0�[����~������G�O������˭��j{�`ޛ6m�O}�S�؊�M�H���/�5�֫LI����AQ��v�9I�p�(t��XY�_�m۶%b<f�"?�0[×V�/�a���
�y"�Zk׬R/��}�<�G��0�U��/.�JoO��-H�|P?7 �]v��e�>7
���`����"����=��K��?�qz��m��>(H��=컀����{v�o���MX�$y�������ꔳ��,�G��ɤ�,��υf�����6m��v�BG���	
F�X�q��iKu��R���]x�
�,[�R�ղ<��ӪaG�qG��!眳M.�����I\.6r��~`߁���|�8����wZ���ɇ��}�p�c�N�ʎ��q���W�'���ty��"��$V~GRg�d�YB�0�o�1[���,77)����8?�/�ɉ�K�������y�1�_�2�JƻX�J��5*  ��P�����Hދ����-$}��o �?&79�lbC�z2T2��gHzs�}!�
��_��s0��k�:�iP�����y�@��-��y�_����~��,��<4�1j�������?o�j�$+d�X��{:dO'��U���Y��(%K���_n�Q�����]O���s�}��������XИp<������=G^�����1Y�t�\z�UF�p���Y��T���˖�%����bIg���m�<t1$k':>������ :,AI����ÇfsQ�Q��h�gjpsb�#?q�����E�M�E��^@;�/k�B+�\�>ԕ��A�4�����m�=(x�~c�R}�/R��^�7=�`ǿ��կ���ߟ��=_1P]s�5r�7&�W���3���]���j�H��e/7K���&,2�DA��%�B�G�߉ޢ^7�F"�}#ȓ�o�9i��+<���$i$�U�A�1^�\_��WY���0#�a��?���������{����<�B��������0���<�ɟ���gC �y���׿���{��{6Ǆ{�a"$���"S�c�y��j�wȗ�����K�AC�=��/|�K���_�x��s�]�?\,��2��Φ��*��k}�s��z�^t�ҥ���yW��e�^���JZ5m���9�Q���6&������-��A�nX��n m�o��o�{����I�+���bwl�Mr7�W����!�[C52�%����䴾[?e�9���6L�h8f�7+}�
A:��Z���(�sB/D?\}�����/]�tV�����ph�ؘ���&�9ر> ��}�I���JdO?l7�kn��|A�>�LY�r��3O�^j��W�=��q?I]26���
E%9�u���S��ӛx"~��38z�b�	;�[�͈���k��<P��MG���,������gϊ�J?,��`�����C�����dQ���k��mF���d��+L�A��=��a�!��q�Fy׻ޕFrmq� �eq����TM���׾��\W�<e�RД��)�G~L����q�d��F�q�� ZP�<ɚ���7�pú��߿�v��B]f͆�=�Ѓ��s�w���L���zF�����#�=jud�%���~�*&
'Z|X���o!�b���UNE ���R�c����p�v�s-~��
����ϰJ���ߧ�dώ!!�W�ӨI�~��' �q8�^�{���`������8Y�ʕ��?/�m������}�[��l����=��a/���'�}eϵOO�k�ϖ덞�=Syvqs���uB@c�RI`��'�y*1�}0�_��,��y�fS~��{;�{ts�X)[A����g��/�����i�珌o������RR���f\!&Ъ��/+V�2W�O,���a�����zUd������M��0�?�iq�9n�W������l's����xa��%c�rȑ��^�|���� ^�������}sh�֧��I5X�xQ�Q��q�p��S�u����a�ؼ����xp����1i_����5���=�䥳Ё��f��rQXO�+9j9�T*�sCh3:o���뇑�^D�P�B���g�Y*.��(� �<BZ���%�^�'~�i�|�s��yŋ���/s�}��)=ey���>ԓ��~����7��]?>��}$b��Pq5+J�#��a�֭r�X请�[�T�ܷ�LV��l��~y����D��Z�I6?�C�NS���rv�:��\�!~%� ���?����d`�	',V$��.C01���OǌX���f��}�!x�,xp����7[�>� ��O@���͍͌P�� �i����`��%�������7==)��5��7�,T
LB#���~7���$)^V^��ot|,��)@1�D#1�!6�zBPњ�9���0mV���9iı��1{:{���B�����Iٹ{�k�L�/|*&��=P�C��8��g�|�)��1��c68'�p��s�����g���3`�����b`?`��0�9�,{V��y=I���مD�yqo����tp���կ�#����~�~G����)-?�Ž�^޵F�x��\j �B�^1�a�����G��R�Щ�:���N��F����?h�v4n�u�k.�6`E�Ʉ.�ѝ�j����|GN��,X�VD�`#�DՇ?�����w��xӛ����̈́�/�N�`;J�#64��f�Xf��惫⸰��=P��l����D���a�;=\6�e2ˍ�����I,��}D��+�(�yh�IbZ��Vz/��1�ZR�^�C�E��XQ��h>��r��C��,P��J��*(N�p�<��,p*�f��?Wț�ea�8yJ�M����� �`��s�;��|��dqds��� ��1���i��� ���F>�=L�����[z>Jέ��TPիr���A�,�$k0N�Cr�5����ú�0/b����"	,�=91e�	���U���I���p�$q�t�I4�ߍ���X�e�2 ��dŊ���Й78ق���k?��w1|8'��ߩ�����r|�()X��_h�j�Э���q+�D���q|��6�����0�ޜ�W����(`}��l��Ij^+Xb-Y7�0�C\�)���{�� �,H��_=���{�Ռ�3gB��������[�:����\�0�G|v\���p�?>>C�|���S�g7/��J��珠��:#E�%�ߢՇ�b-�o �d2j,�l����&��8�,e�dB��ϲ���{b#h��u��ۨ���?V	�^d}1�0m�� �;Xh�]�X�hcc="��x�ܳ��f�=��C�@�x�Y� a�pQ�R���̑l~q/��(nf��Ru�h?��j�q�)���KH��Й�}V���%��;@ZY�R7��������˾��i��L濓�ϴ9tJ&�vt a������)<�P�<5�����o?gp`�#Wt��Xx�� �\g&��D0֜����3	�3p�����Hl�ÿ*?�M���8����l:cs��17��ʦ�4�e
�,��!�Ű�M|���,�<�߮/�p�=��a�{°�	�<�.����u��3���	�`��&��ǉ\�9|�;�� TuA�Z]zR���w��m�W�@�$��� 7��o�/}�K�w�ð���c0��_���>��ǥ�ǩ=�}�C��
a[`�ִ�o�qӷ��~��k4b���t�7�ik×ʹ�?�8兿�C�0s2�sq������`��ۿ�[��9����p��C�dl�H��!������g{L�F�
lME���j�z�=~�G��>L�'w�3LO���A�������� �+fr�
�f����9�F��D�I�8����6��)0��1<?��G��虑	����d����(L�g}�b�q���sz;�<��6�����Cs���������W���y��<������V$�O�q�8�HY�|O�3 Ny��A}<�`6������b?�O4F3���P���ΰ6B�D�l5���������`��,n��(\�h�}�͖}̤S��1�n�3n<s^�1��;!���Oo��'�s{�c��ii`�u����`}m��Ux'#r�ۢ�+��)�g.|���'�����M�4��h	�0�w��k�w�l��~� 
��
^
@=�io��s`���"�t��|@{�,��Ѭ����_���?}���Ж�-�F�	|�ٺjSP�{|�%ףUT(�ݻ�����B�R=�P����B|�,��9}�d��s�܍ފO[܌��B��z����MFG�J'��Dn�|�x^=(V�2\f?��̦������|�����x�,��I�XC�b~�c6�?9JGR�T+�����������r����>�oQ��lI�l�7\�1L��I~ ���Jȟ�E YR+!�$� �)�1`\0`\�1��]�,ٖUn�w���g��9����;�;��+m��\͜9�-��gW5�?���U+���bZfO�*`A�Ey����.1�l����[)��a�;�l�5�GaY���H(���cQ��p<�-���k��7����Y��{�ޅǰ�����"�{��P�4�y{^[�w�1~�����W� Vڣ�#�}c�+m���?��UuN�W��ZE*e�|Qq�^�-�w��m
c̊;l �����+�u'j����2y��؊S��Y�ąN�*�����8
��Mt?!c��D*d%�ez`�<m��1X� e��8�}[������0Xm��%K�m�p�Z���,��D�sT�����sl�$���.F�<�
���3�56Z��(bKgRzL�Z� ���#�(1p����JX�F�A!Bs��.P�Z�� � ����Fh�ز�N�b�(qL�R�1�B���9f%lR�v����G��9�t�b,��7���x�	���8�}.��sj���ϙ3[Fǆ��zp���A�]~��q��ߢ|�VK��!�дg�A�WD۱�0Y���}�\v��N���Z.)�b	Mݻ
�Ig����uN  �1 @�l��
^�fc!��Z��GX�YL��Iu�����&��N�Q4�U`0��Lm��u,d��dT 2A�q`�)Y�KfNm�V���"��Mgb�:��Η��,��d��r�S��N�	��1��2��Z"���ñ}�5�Ԃ9~�'��ٓ�<�!S�q*
y
��5Pج¦���R����� ����պyO[0�}��h�A�ь� pOj��5HAa�/�OXw���7�Y�
>��,=�9�u.���Y��sf͒׾�5���\���^a���S~6��4I�Ƅ`�g��`yL֟z���Ȭ�3�f������=�ec1\��c����9�Md�6ky���._���b$E��� �a���B�Z�&��D�$�؁��K����d5C
4ݘn��Y'c�8�#0�!5yj�d�8?z�W)Y�O��M�sw��59���ٳba���иy��[�%
�;�.BQg�g��92�����b�3\PL ��X`�cQ� r� b�>�bT���xˠ^-�������G�f"K�L������L�������a��D���&������cl�P"�Nz_�����t����]�O�tQ9!��U���_�����%�8��ݷ�٧䷿�[��t캻���h�)9��c��7��u��k~$/�� �@z��ml�i��C	�z�8y̓/<_�͟-��N����~%[�>+%'�!e+���9&O<&3,ǝx�t��ҎPhG�~lR�?��]�SN9E���_�m�K퉌����$���"2C0	t.BĶ\�ϟ�-�;p΁e4ٽS_�j�\v�eu�t&��Ʉ�&��ǀ fs�A-���.���Q�̟Z�O~z�jRV3�1�
�L�-'ў�`iDs%�0 ��o�a��Dc�p�b}��K���.���C(�X4����C��U���M
e��s�9G�=(ȒZ?^�=p��z��x���S�Źѥ�!a�R8[��>>��kY��f�{B;�3�<ӯ�Tz�rD`3��%q�/c�A��ޤq.4�w���O��|`\<Hm ~���uD�� @;̕+�;!^t��O6��<������(� �z��k�rB����M���;������B��`��� ��YS�  �A�-���\9�%R���}���e��s�;����-�����'w�u�l~�Ey�;߫Z��@�>9�(�t�^{��7����_�z�h�� ��_�<�7�abc�'�	'�0�1�Uc5i=4<S�����8���<�+
�]n�yO��غ	B�q�ʬ���jo��0�?���4��P�h�y�\U�����f�02+�0&`Rt���E{>�#�9s��r��hL���)v�^�����}�m��*��i|=���cM���E;�ItS]�c>)�gŊq۴�������Bj7#��&�׮�S�y��C��82ִ�]?6 ͽO��Z����ZQ{��1f����G�޾��o�J	��P��k�S �,�?z�<��S��9�;��~��<������ʍwEN[�T���=�|y���Um�|L{�6���is���渍}�G�s��;n�#W-��;�ir�ed�_��7�G�B�� �<ޠR��6���>L:�p`� &�@7h�hm���7�u ��6֯����t�n�6H���b�H�9��[_2!0o��Q���vM�ic�Wۀ4�),,tv�����b_./]td�60=Q6�2dtn��|]O���0%�źk+_p>WPE��@ 
��1j���0F��gLJ��͞�-3�5�y�:����S+�A�ҹ���x�Y2ѵ�?�k�
,�Mco�8�vp�úB������WW0�� ���|򓟔[n�E;�q��~a=�=��?%�g��Z(7=	�(�+ȩ�Y����W;
._v�
�#�X#����[;�)W�N{��,ϟ�L��×����twed�K/ʑ+�Ȍޜ̘�U(]��LAd�Z��c�ve��21��܅	�f4�|���Lr��.��b5��XsP+AýMt=�O�m8������l���7HR�M4�z
�����Z��q]��O����y-�O�I��P�4ux�
f��x2Qjy4�q��lf��d��k``� ��x-��6�)�`��ٜf8"�}#�$÷)�d�xv4Ɂ&��r���B�)����^���Q�̙׎!���ϛ�}p�����Mg���|�l�5쫽�?x~�g� pK�.U��������Ö���B�p(��7��`�6�>"�g�d���2w�wÏ�X�hA�����-ȝ��[/\!�3g����e�aK���Ti�3�f�����F��;G%l��-۶=�-HA;F�v�;I���[yL�|�8�S�`�Ϛ�AƑꈺ
�����_�1����Њ��翐����̙77�Y??Lln��I4��t�������y�|��Ǖ�=&���s�E���q`�b����:'s�)�d��]�
�����X��6��f3ڋᩧ���$�;�L��ܺZ@����70(���������3 ��
w�r���)�C!±��êD��fy��6&���঺t�z���?�-/k�P3��q��d����a�ARY�.*úRk���M�m��b>���*��C��MoR�/�� ı  ��s���^{񅗜U��?�(�g���NȎ��q�"�q�Y��ky����.�M�����_|�y�Vp����h�3�Qbb�v�ʦs��Ckԁ��lJ��ɡ��c�5�ӒqǏ�n���Q�ƄM�F�^2w6��d��M�l�9��=a�a<�,��5*���V����O�qܬ`�}um:� �^��8��Ա���}c������cj���6va��Y"w,	0�fy�,X��F�<��gצe����%ƿ'"��®++���I����"�f�q��ʰnЫ�3���|�󟏳�p����ަ�~�/��8]'N��#w!Z6VkN�G6W&���J��`�qp��)�t2���5�6':b<��O��B
d�8�ȫ^v�
��g^�Їv��wҵK���ag��iSK��;�ͬ�X��p饗j�j��@0��{�y�7d�gf�X_��$n4�dL����J܂�%6�f7>c��L���[�i}��\N �1�c5P�l=)sh���8�3�+��
U��-�i�67����%%�k����c��4c�v�9�|>S2Pm����#�wؾ���xnd���_��j��v���������g?��c|i�0#��B����3*�rF{���ު��yi�Q�@]�iY��-�Ҡ����S"kHR�0Г������x���	�_��	�/=��=g�̞��i�nӧ
jrժ6 ��K���\�Grd�5�ό�{�G}��}�k��;�6rva~�+_����7�f�Y�n�6���Zs���u�-cO.�F�d5�fZ0�ϑ<�-@%���Lx�d�Q+4��B�g5|^�~�8s�h�Xo2��˞�ײ��^׎�i(�~3�k����K�}����J���L�eb���e@7yO��ܛ�k��`V���뿎�'�� Ա�Y���cb�
�×.��b5-�l |"B5��I�`����󥧷�E�>�E�B��[+��q���?&o��5_������3ϐ�;v9F}���}��9)�#�fuG�+9YԻ��Ԟ�.+V���-$9Z5R+����P� r�!>����>�1�җ��ھ�ٸ� h�l�7�'%�o�_��%��̈́�ua�sY��M��Y��t3q��2jF�1w���|�y�6Va��V�?��y�ɿ��������
�f�׎5��H��9��[?=�����co�CA`c1��j���]�E��MaGK ��9���{����p�����@	��dՑ�ep�%���B�L�vVB��U�Y9��3���k6�G�@�>�X���$޳�0L��P�����\Z�{��.7��{�L5ǰ��966$4fϤ��v��r��r9�����0�M�6�@N�h,��.�*`��?���p̒a�������,m'�!��Z�e ����2U�:HZ�>�L�j��Ѫ�Ԉ�l�E���&�߼n+���&yV��3
C+x,��cb�Jj�,���P�ot�V,��{.�Z�1Ѽ�m���B���(vC��;3߬0~�ޠAw�&p,���:J��,;���T�Y�R)�M�1�h2�ͻs�e�;�s�tǮRK ���[�QQ�k��:o�WUZ��r��r�mw�+/8_F�Z�d���"�������c
]r�I���^"s�-t����wOp���_���wj��~�� @̶m�����l}���bd���w�/�9��i�$����ؤ�8Y�����h�[ �%��O���ǤO�5b����`�2+k�7Ҿ[y������3��cac��ڠ�T�2�F�9?�ț�[]TlƘe�������v-���������KZ�M�EV,y$s�uI%�{��塇�SO^'��,9��N����]���������b�r�y���k��r1����]�=*]��b�Dn����?�?I~� �'��?��P��c�s_����\�������ŭn�f���9��8�U��� ����=�,���0�9|���*�׮Q낛�n �q�O"^�D���Í�{�I�}���=�s翭��U��H�p�m�)���p{��>R��粩�I����
~N렙�k�u[��<&7�s�T�Ɉ�g�xr�W���Z���fa �?��?W�>g��f�� H��;{��\�J
�9��3�UGɖ�7��� %��L֬^�, �SR9�%��#���?�ŝ5.��s��V��=�oF~��9L��\u��w�Z��	��9G�Ξ[߬nB�ق���u�}/�������?��?>G�=��ƍ��͛b�.d���.Y읤o�L���`l�2�F ɸ,�� �����>P#�ОR��Z�7I�����ͮm�C��7���jF��1�&��~��o����a�k�m��k� �}?p�Dw�2��ـ�����A��
O�������7�M?��gH�[����I'�.���xP�]#x�P��n����:+�?��� ���S|�����^�.`g#0s�q�)�6�}L$.��6l�GyL�=�0���l,�w��ݺP�@��8��?��'�.�={v�;5�v��� �8#i�X�8��QV�>D��`%�ka��}ٲe��|�f=��E]$?���!�ҽ����{?��b;�q��b�
�'2��/bk
(N���=���Nhx��g*�B�z�N@���u�W� S�7C�vI��}� ���u� (��[�@ ��>@j 4���|�Wj��Ƣ @�> �z�ߨ��XP� Y'���
�/Ns���Q0j �vb�:�S�a�#U�C��Z�@�E��x�`�Ŷ��a�Ê��������C? �;aR�g�2�*j�V��R�r�_����ө��N�N���G0�Aq�"Xa���&
�
�Dj*�7Z�����& x!ЋB.��~�a�馛tB�����f! �:�����Ad�eQH�F������Ƈ��Ob�������ܢf�+����˿T�
�u���� �l����3}'����ξ�}o��4SWÈ��aӞ�7���<`pA, �xV2ٌ]@�����t2Ku@+[}���h�$����=����;��&�M[#=��"3�=D��`%��2�M��1����������` ,	��{M�E+�?���� �֮�����[��gS�q�FA:OL�g��|�8�!���Zq���.��-�3+�S6�[ڝe�������XT>@�"�EĎJ6ۢĸ�f��%����{��E~���v��!���p�0����}�s d3�\�f��dVF*^ڗ��BOlex�>�k����PZٞm�g3�OGn'���R� oZ{�z�|��K�4���E��v���_�O�ӊ� ��XLHE��׾��* �o���ЮۅZ?�6����l6������=n�OX��`05||��O�~��/����f��|�+V|L�1`��
�y�@N�{��LZ����'���D�i�	���g�M�����]��N@*=��"�Whְ�̜Z�L>�����҂�}���"J���4PJ�$FK�f~�h��)��ŋ��� �������E�<���5�O�8hNcކ��ֻ�Ѻk��`������ҩП����/�l���m	2��=��f�Y�E�3�#�^����7[�kB�q��>��<]�A��{K=B��/��h�	�+�@�J=��~�z*�׺�ƶRZ�D�02��@<V��oP� 0bҷ�ܡ�$ѯ�ģ�3���(��^s��=C�;�X��e�M|*���y�X���cŇ���@d�X��Np�=�j��e�,�T}+?x>�r����z�����β��J���촞,Vp0E��^)'L��3��� ���ZM��N� �k�]�ijn��1����� ���[�)����U�xR���@�琡ں�d�� (�$Pf�AV�K֊���bƎu��,�m��?����[z��]��]�"~�N��sLg�S�����L��aJ�����[�!�hzІES�g	�,w��ò� N��G�x�z�"��Mz�p��DGc�^K��s�0��շ�yj�48'�o�vl�
ٜf̔��fh�K�k��cJ�RHd��E�ð���;GB'�*��ҹ,L7񚿿�={G+Č�`�Kѽ�:�e�J9�-��0�}G�����/�K�_���71H��t+�Aºd&W���@!�%P���s����O�Ly<{e`�����R3EN[�"#d�5~>�,j�_���ղ��T�h%���󟴁�����5�)*W�:I�5`/GЭ�jݯO���:�m��V�"s�����M�DR����A����YRp�*�����O#�F�;����>;%i����;�̌��B�t���<t�8�T�u�A�,��|���쳲t�ar�y��9�,����NP k
̿
�B�1�ZQ��[u���-U�W���H:�J_��|Ӎ
ّΠ�O&������q½w�*�8>��F�,5��}E�_0[Z�!�M��(`�x�����T�|�[8��dd-�F�t+�L ���5x�*nQ�O�[�,�EJh���i��C	�b$@���ה�����3#n��H��V5���v�I?i^'K��6ɓ�k~x�Ө�ҋ����n0f��i/�]�E�Z��eo�_J��ݲ`�|��;�i@�R-"���4�XK2�Ǚ��;�4�Tg������E(�� ~��3�����	*���䶕���fc�nӹ�̘�#��,�o��Kp;���@�FF��B��2P$0~:P\=�p���&�L L�%���SH4�R?�J�e���GX�z���zu�R�F��z�(�<nw�Z��k�!Ϳ!�}zٰ�1�rMq�1��C�n�u�.����(���}n���wO]���mTQLַc�{Β�YrQ�?�}�i��%g�h�Ϩti�W�� ��,�h��~{�/��Iw���Ԫ���^ɧ�B�He~xǂk���!��.�9&0�"NVkS����g�?W-�� ��T:$�ZY��9uE�
y	�Z��Q�����"�XM�ʽ8U���Gx�LCf=�Ex%fՁ^����
�6k���Z]�&C�X��w�8X�*��4Ѱ��������5p��A�=4|,("+
����n��w�1�Ë��M�����	[���b2�}���G�9F̐l�G��Uefź�5W��xn��3��*B�^Vj�蕙s�h���`���%�<:be�7���9���gܳ�z�%ǐSmdD��i���ԱgYcN<S�FS���	�J�397�9't2��S�b���|�ΠӚc��D���0�FOk���`�׶4���E~�Sr�'�1��؈,�?_+���fb\��B�W����6�ӰKQK�\1�������>�h��[�MY�l(�)��ŗ�RN?�tQ=0J���>�9�u���jr{ٮD�dU��Pۣ���Į5.�ae����$К��������1�*�����o4����vz���hmX�8m>���T��y��s�Nh�Kge�1�.�}%�I&�չ��v	�4CrZߝ���
��sK�{�.'�rRvB�\)�X��!˖.�MO?�kb;4I�4����9�:P�%d�̘�#�'.�Ŝ�3ئ�:5�3β>��3��sϓ�n]A1�
�`~u��ZIL�������}M{���3hJ�ޞ�����sΕ׿�5Z�U.�jZ$�%�"r!k� Z��|��_��6m�tO[���i�j���+9F��c����qV����U  �"�;E��ct%�}���p#�qi�PkN�h��H���tI՜�VH���G�2V��ʘT���v�;�0�B��˘ȔR=5[��-Q�eU�⳺$����L*�Wh�1��~֢� 1,�c�����u2 69gS�|�Q��ýv �Dֿ�72Yy��ީ�������ݏ������w) ��UGʯ�k��m��|��.���D_L{���(f��)��"W��M�Q:��M�T�n���"}�}�`��Ys��Xy��dg�q����ۿ�[\-�I�$����?��?��~���'�&�ැ�>L՛����3L�Q����n仫pH��X�� ���{ѣM�8�B������$,�J�����R�8�;�>K�J-3&Eg%Hۚ��}G_�'�jydB��H�+�Vk("s>@�T�9�WM��+O�������5P��n�U{y�`2c��݊{���P�t��u��l�e�{��J{'��I��� ��Ś�~���mJ�e K�{�ʕ-��P�9�����K��a�ڬ?޳���1�������6Y�z� ]�/tV�}�<�ݼ0.,�#�X��u؍UY���Μ��f�k�<2�n�3��ɾ��x��*K�,��^y�t�s2sV�lټQ~�>y����o��Du��'�g��Qǜ �ן����e�]����s�9��կ�a�� ~�t��o�]���oi�7��Y"֠��h�M�{J��:t�F�J��8���0�i��U�V�-�·��L@�&�]x���>�.�2��Z �4�`Yw���G�1��%���R��ߖi��Z����tYw�M��.ٚ3�L�%�J>�M�`�<S-z&]BG��Y+�b�St"���H�<@� �
{�9�����p��_�=�0 �/��r9�5Z̈ڢMO>��Z��9�:�v�nY�r��~�ٲ�5�,��;Y1�  l��Tb�Ӟ�7#g89�c�`h����Ҷg���[��#����h��Ӣ�����V����}�yH=��3�_ߩ�`,
hӐ�-^"7�|�B�b°@������=��3yV�/j+,m�7�Oj&)��\��(�pZc>�6t5#���K���s�������ˏW&���VI;��7橥*�ʨ� ����^��� ��J�$�6��d۞��m�62(��j{�&�M�&���70��ɸ�M���?�LP��ReS[=K8�N=C������rꩧꞇ���/��b�����=�ZE�ݬ8��ի���O�տ�rܼ�Qyⱇ����+�?,�-c�J�������ΖSן�	
�7>����r��^'t!�)��g�M*|�Y��*U��a��淿��yY�l������^ �<�B�ᑊ�x��r�jY�x�Jx4kA��>K,��[��Yg����������?_@<�І����tM��{*�aG�Qq��|v�P���@Z�5rbld؍u��AT�&��K�?��?A2�j�pM�R�Z��u��b����1�q�5W��ـ!u��+�Ȃ'2���2:��0%�{��G�s[�oߩ�C�c�ȯ�JH�H���%3��;:�&�e1ЦA����*~��R;�1J�C|�d��?^>��O��c���Au����~m����^}�,�x�*�]��2&�f܊*h��wUah���䦛n��K����T�@�`~[p���nA�?'���eK5�6�Ч�yR֟r��.[�̲�8������;�\�J���>���;��|�n:�k�qD��"��w���՗�n��F] X�X�����$�)n{N�l"��tE0�6N �̘׿�m��RM�-��*�28�]
��#�$��|4�ew*]S=� R1��B�3��0��V��!H��ޅ�S=}͇w�x! �P�RtLi�c#���ޤ$���j�I'��4A���?'�4�� �P����:��q~��~}>�ʗu[��x����b�Y1�2|@r���2]tP����	���к�u�E�{� ����/|�ʨ�	H���ʕ��yxý�d�Y�h�����;.М�+����s,�����j�W_�Z=Ǌ+���v��V�m�3�fD�����ӧ����s2:��&bT*U=e�\q&fyX���� }+����I��,6Ӯ]�T@@; ��{��^��0�&:����l�@�|e�@�t&u��$Ԕk1��~���'^>�rԴQN�<&)7���ՃYb��`��s�"��? ���PqO�ӵH��"�Зz`�0���T �� i�C��F.�0�Ɉ��9�8K4ɉ����,�KNͺZ?��.i��F)d� �8X�\�{ҵ���<7����ۥd�&�O���x(rK�.�7���կ~5{Z`���Ν?~�ȥ��m��='�4�n��lA^�a@�c:�1}��}�=���/����W;�0,���k�Z Ӟ�������g�%cVq�3jv��	(9T�l�riDjUg�� �3�j-@*��ɬ��^��T쟋��O�S�����MDs��K����[9t}�"���BA�cHtu��m"�����h���͂^
�ﯦ�W��UV<� 5����%��DA�v����Dh��T�sBp�v�g�����^@���MnR[	�,��-n<�%�y��$��[�&�̶K�G�;��y߼w
�����a,��If�gc}���+�}�ϡн�oTW.��ڵk����C'�w�Ճs ����~��R��}NX��Kh�@JQu5�ᾃ5��R��c��S��i���5sa.1����TN�xs���������� �����G�)Mgh�0����oD���h��Hjm�ק/�M�1�8��h?��f��>7_ǄC���Hۍr�c5���5��w�g.�CuL����!��(����
����gS#��S�o���#_��Pg)�4�S��8rt�(�ã
+h�M�L-�W�g���p5�����M��mj��NQ����Z6+Ǧ�RC��kƽ�p��a�C�>�ǴK6k�����L���%��O��
=���NS����}M� ��e�ݧf���W�������og+I�si�	�2:6,3zg9!��1Z��JM� O{�N���4��]2:R��+��KfΆy��4�R)#]��NW4ҷ��Ȁ/RM��/���1�!��W�*2!R:i���X�h�UW�}�&�d�%�.�OM�����2���̛�)դ�������	c�"恳��+ձ��s"�240���,p� ��F-�� �vL����W��uB�-���5�SH`��J��[T�@� X.元fi�����r26<�n������QAd���t��y�Mx0Ƥ4VԂ!
u��y���� ����|���V��H �:�<���$�BbO	���^�����تZ���x+��o�E�������[������;]W�����E�:�(�\a�޿��䆛n��R�6��4Ȏ];=�������e��Ŏo8K��B�L�o�ҘS��&�/�X�ם�>��%�Ok��j>{B��BӞ����cOl��O<N�֟z����K��]n8!���M�O�����)�y�n9��T���7���>�nL2���ju��
>Z�數Mls�4��B0��dұ�b��N�F�r�i,��1~�؛׮�;7�_�j3��+��(4m�<���������x�1�Z��,��9�|V�n�T��L!�'��Ouų(J(�Jj�D�%��1�����J��r���u�:DQi�Ϟ>|*rxG �>�|��?u���آ��B7���;S�=�x)�������~�2k�B�(��E�9�,��v�ˮ�a9��ӥ��[�d[�<-�7=%��yiFmߠi�bM��0�P�q������Wʖ�7��%-ꁦ72:��9�[4K�=cr����J\,��^zI6m��4�L���ze���C�c �yx�[���e��D�����[<���F͛+����is�7	�-��)t�E널�H�<���x���b���{��k��KP� �Xq�1Y'ra�Z�g'�Tݴ �\r��C.���X4FS��f,�mړw`Uſ����ܠL��-tfKe|��������b
^
�hjd��<�%Ō=ya@!���lJC��'?����}�,=l�<�н���!w��S��d��T�Ȃ�K�R�ʪU���/W�cht@�{�Y����'�i���������=�������'+^�����A��'?���~�+SJer�x���կ�E��Љ�tG�|�4�p�򗿬���1����?�o8G3��

ݲn�:y�Wz�(���3����w�� ��K;w�=�/�n�VՔ���)�zqc��-�1�7`�1e��%U ���6�H�1��z���l�dr�,��F�v�m�]�WoF{�jm�"z[�YhX5�a�k�E���;����d���3&�̝׿��qj7>g2�7��͚��{�Bb�ƍHϟ��.9��u�םr�-�r
�f�UK�\�]
/���s�=�Y�0Y3���Ɇh�QOWs�"���_�d���85nH��{�1NS^�����i�ٴy�j�k�>F�S�1{�cZN#t��-��"w�u�8�%,x��(?\<G}��@�lذA#�H�1V1��%����u�a�d8Y63�L��E����X^1���%$������w&�3�Vא
M=�ˠV���/�Ɯ��%��,��ze�PU������vR)�j�=R^�=�ŷ���yki���K p�iphX7�:��(7]�t&j���U�}�L?��u�?2�Ps��B���ه�d��{�ys溭�-��~��Y}�<�Ѓ�e���e4&�~�z'4f��pEQ�~�Q���~���.�ixƔ�M�;5i�D��	#��������G����n�3w�6MX�t��x���#%�Q��M7��Y���?��?V�����r饗*x2���
�Bї�a����k��ry>�b�����#��p�t��h���6�{ob%��묍�'}�04l�!��2&��(/>����%ya��̎T�U�3�xr���'��3�>�<';�������0S��rJJ��t���������MU*v/�C�&Y�$f ����Q�����5�X �:R������D�R��P�|���hm��×鱳fg�.��pX[8N��s�	���Oʏ�cy��-*l�u�����R=	�06R��z�t}�Qg;M��x≲b�2͂A:&�VKI�1�ǞxLn��V7)��0Y���DÒx�k^����|��؝��я~����.�H���!@��Ru���j�2�L./�<��|��߈����,��b)����3d=�:X5"NۥޞY280"w��^M�����ל�)���$�	��������f����K*�U��x
�?��<�V���w� + Up�A��|Je:�#a��Y6�-�h��m.c���R�h� w��m��;��"�}�yp��0�];�� �p���9��p���(bo�xޝ�~��/�����V�i�3�s���B��]�9�����a�͘5S-X(���v3�]��eǎ��s�7��n�219�D�Ϣ�|`��|,X��H�p�$�7p=Y�f��C�=��(\��	��)bQD��!M�+��^�i�t̠���z6ױ`����Yݕ�\
n����K*'�3��҇�/�dj2�/�
|�.oqQw�s�V�*�=�1�uTS
5S*Pl��gZ-y����>�O~��'��Q�뭷j���ɟ�7����"o�;�Lxf�32tː
�U�V�+�T�`�=�͛6�s��
��JeU��+|a_s~�������QGZ�x�	>$F�ˣ����;�駟�A=)����Ro���(s{Y�?�����%D�V���3�tG�ԑ�j:b����ݡ��s���q4{:=��u*�����4+Q�^��, �U!��u�⎫��X�`�)�RZ���L{��)���x�P-B_��Zw\{a�{\CP$�V�����i�v2-��
�\��tF`3n�v�&.�)�դ[ (��<?�W,�u�r�9x1�����~��T�����;��P�
�7�7
���}H���'u�m�7!]����e�6 ;�v(N���(�5֨�)�u��Ti�R�
��ct���2�[��3|b�KVPE���.0,>�>�я*C�������MM?�zDqd�"��Ͷ��m�����	���)��5�`�&�mj����}��
��_�����>���e�M@���C1W��+��̰V����;0+2D
������(�m�ʒhU�ձ�x�,f����$i2&N�TiV��Q����;�
|�����a��YP������K����BRp�"	�Z�/x��ʑ���u���ǫZ���p�=�oV����2e���#�1�1'��X���7n� �,lD,@��p��#$�+H�0գ��(��[�����ׯ��E0��[�'�֩E�X~c� Ўc�k��{*J�4g���Ƨ��Z�lJV�-?��#d��B������g��WŦ��*�����ݽ*[�`tP|��`��[�S3�ռ���4{@TX�v�=5��A�'�GsX���D� �{��+��)�Uů皏B�.���f#�i���u��g�惻�o<%M�o~���S߱���ޠ��WH�[|�����ˊT����R��~���?92a�����7��.�`7��CVӷ���$Qx�+ΕE��-*�?RG�"��K��G,j͚5��!��$ԠS�:g�&���I'�$K�,��<�ξ]z�]���F�3�=n��A������(�!g����y����{$v����kt�ӕf�(���\�!�P�nӑ���h؉�9�s2���qI~�1d�5TZ)�̮`�O�'h��8���K�����e�Ų�[c��/S&���b��[^����Jf��9\���1�w��}}����x���'1��Jd��] M����?�~Z����&�?iER��4U� ��?��UK%�&�'R}� �糀�����8���?1q��j9��3�x��`m�r����JVp�E�s" ���~V <|��u?P�������O����_��3И��5�-�	9��g���.����C��lAl���0�B,\ &���R��o�y��q�Zf�� ������1ל|��˞�:$���#�v�
���h��&/���od�=���2�aЗ!�HZ�E� ��v�*כ�[�xOt�C�h-
4SɁ��"d��פ�<Y���q�����cQG��e���n�p�?;��x�y�6���.� S�����/L�s&�SS�i�������:9�c�o���8��͟�b !(f���\b}pS��	;aj7�ĭ#Y�x���,�i#��=�8k���� f<@�bQ'��*���@{�>�V��z������RKK��o�
١�B����z\�`��7x4�kLW�:�dĠT��ֱ��!�ݟ|�ɒ&c��;��,$4�k�'
��-Ȅr���wr�;����O� �j�������>�A��7�U2��2a��%5������.K� QK�o!�9�,*�ֱ{O�ERs��x#�_�f��e��߇l��g�}���ek�a܆i�w�駱�t�A�̔?x3  ��IDAT�^b��YٴL2
�yR�d�N:;��e��K�Rq�!2ie��t��h;tY�	�;����e��{A��B�;��ĽMal����g�F��_��EAPW�gQ�2�%��w��V|��hL{�?��'��(%w���b��	Q.U�HWf�T��er��q���S�b���Q۲B�fh�o��-)�*���2��)u�XF=�9��ŜC1�=dD��itD�*�cΧ5O	�^����5�r
!�J���w-ܝ�m����):^�Y��Vp6Ef�6��rkѻ$�Sѻ��lΤ��9�c�y�f���oM*(��1?2,e2)_���	+�5��;\3͘';e1œ~ ���uL���je|FQ��3
N��P-���F�* ����;����K����ɂ�L���+�?,]C��	���e�<V���A)� ��|�7�r|A*���3~�<�fn���$b~���Iiyu�7�@g��bE+q��2����hS�#�[m��G�Ķ����ٱ�������?������}t��� 
�f,)�fY�(�R��|j�A�B�C
̠�3kQF�z.�&��B���|�)�L��g�5{����m=L&?66o\\{FO�2�z���H�g��}���̦Y@6�+LE�ء�Z�z��`�z�S�����l�;d�螱��{�8��Ne��:���;�7v��9IE-3٨[w</P6�b���B9T�#V�/m[.M�ާ=�o��s���DE�:��A#�#��/>L����64]wf]��m?�mMlLl�v&�mۙ�v&�m��}�u��9g��]�]]���[g�֨ ���p�Z�+(i���Tߖȥ G�M�qdM��2�0'��^:x7-��R�af$eS�[���"*D_٢U����	�&uj9ad-Gv%N(BJ�J����
�ǎ��B�wh[��zZ'.u	3��c$��6:qd�l��&�%�#^��V�z��˚93�ٷ���g��Sq|ܥ	���ʦ�&�8Iz-/@<2��TG���<�߬[��X�j�jZ��U�������q~y�J4C��h��"]�j����R{rU�R��4ǣ����T��9��w�Ļ��<q�;�F^���.������LT�"� =����<4ƙ��+�����"�+1�>��T��$-�*��y�D5Vr�{�l�:�r�Ԋ±�Ey&�����1��d� u���b>�ѐ�N/�7AaU��R��o�tY1�7㻇X���pNcf�Ov>6��þ�p��wH�\��lI�`��I4�+�=�J��!p���s��ɰ�F��X8E�8�SԞ0o3Ĳ;(�w$�J�0�'�%v���
������ 9�:Lf�Wew���c)����p�"Ϟ�Ê����Xag�5&A�H�� !O=,��{�s�Лπ��.�ga#6�J�	���������-�%qH>Z���ϗ0_rP���R��٣�!��H�֛�P�E���7>�ic�����v��:w�:�I$W�kj�o�*w�[vq{��ͼDM(��ʗy(�S�}.�AO�?�p�����i2 X��MB`<���P9:�1o�}0h����6wp �4�\t]Q��@
&uUS:F��f�fD�*��y��Q�y�kSnq_�W$p�^�����Q��R����^�_�<q_�e�}�B	���N�o[3��!#b��V��.�e���	�Ȋ����~��e.�a$�j�\k�����l:�a�K�8���d�X��y��e���s���	$X��D����Y��S���p�?��B�i�)��F���Y�*
P`:RQh���e>��!�mN8�Ev��q��B6�~#����3�-F��������2�������ҟ� �R��U^��~�+�^?p�������濑B�����ݗ��o˂Y�Ws.a�J�b�Q�hT��'�]��M36�U��4C�'G���{wj��r��F���!`u����y��)U���>�a;����f#���UԚ�H6�뎛*S%�;ڼ<��3�Y<K�6��������C򬷟���d�=w͌�c����b��e��q�(_��1'@'>+�>�]�@���m2�ΜY���c*�x�z��T�S嘎���Me���Od��3ǔ���˭:h�l��1O�k%��S�:��쬧��SZ�ݾ�]?����S�ܽ�E�/�	�\4�M1��6_y���d�j���Ue1���ѐ��Z���,�j+b�4W��d�aɞ���D�����qAL\K��_@�q���s��Zn02��k�4�\�k��<6̵���[+&�$� �>���k�������� wf�:�V��>\�e���x�����*�;�M����F��g��K��;Lyk�����Fe+� 5iQ��.����4�������/1����Yj�4n*�����u*�֐��P�ɿ����w{�����ϒiF�7?=�h��.�bW:��Z��.�� ��U���ˬ1�x����Y���Ԣ
�W�ߤzB=Y�B�^_{��9|vڤ���%LuyU�e �-r��Jڷ���n����(�8��rk6��q�Aec�\�L���o�*��DP�m&O{y۹�o����8�3���Bi�H�~��P9�������/�*����3�%�#nR��ViӞ^0g�>D��,e�T�}�:�9�i,&y2��^�8x�d���4U�pQ�0��8a}�K��``������F[�2c�K�QW�n?���9�>�~?��nkw��-��������}_��}�8>�i���J�� +��L�=c
�+�X �kdw�4-�
ʘ��9I�b?F&�s��ל��本�">�IoL检�*Q�[|�ɖ����c����8�&,G��d�}wJ5
	;�#���q��t�� ��{�P��w�-a澜U�� ��@	���?z�˸KN�|�}���͜VK_�Q���?����ZE��~��}�6[���f�f��ߟ��U��0Wv���c��Ev��Q�	�YH�"�W&�W�B�xc�����RkV5�-��x���������z͊9[w�<����e�|Pi���R�<��q*�,p��*6�n������&��R��q�
�v�s�z�q��=�Uv��u��\�'�������i�H@7���I����ӱR�V�֋���q�$�+�Sw98H�t"�y���ݳ�|�@�ٴ�p�+Ŗ���P���u�m������Xzl���Jp�� ��B�m���=%����:��"������&k,4�}c��I KW���Y1�dx�O�ϓ��zM�>�zUn�Hv��/x�6�XE��S9�	O,�����PP"��i���(BZH�]l�n�"�Pnr0�i���b�o��$�Ѡ�j�Q���T��.��Ѵm�~�1>E��浱se�2^��$��w1��P�h2�Dt�oh6y��:ltL�3}P��<2����t�	�/��N�(��#x�bL�����Q��?0RI~U��?&[g�3A�� �M_F�I}7F���}a�A[m�/���ؠ�p��o�qD6-"'�_��t�_O�ze��sT�妅�t[ބ���؂v��~`��Pq�)�)��&�鄲�~�2-5ڐ�# ߫�D[��QH0�P��e~�Vy�I��C-�L��Lnk�6�a��s�7��}օX3o���b>UY�3}ف�u��ߟ�V� ްU{���@w���C�t��t^��w�*�gH���Y{iǑ0�\��~X��6�:��!�_6[�Օ3<'lߌ��>���'X�&Yy�4xOʕ�5�M�iDc���`���k�`�0qA	�7 ����I0@��w@@���'3��: �D��q6Ap��uX��R,�7qş� �N�����9{	#v$)�8���Z*��s� �������=�[�9�[yK/]���ZI����.D�܂K6�M3��,��r��G�X@lv]��.˹]f�S��T��,E�pQxོ͕K�m�'o�;7��\�1!2z_w�lN��������� ��&����v[�a����Ƀ��
�d��-J�����,�vUP�?�Av'���/-S0d�����l�2K�A�ړ���u�N�咕���N(����j]���O+"٧6�<�O�7��$ޝ���L���,^!=60��E�9��}���agM��%�O�4���b�ˁ�^b�H�{
P눻�#����v>iX3��#W�^3�_I��r���I�6�lc�����p��n�2��v�����4(i�n�d�N�ˢ�3ރ��+���Ӏ��řp.p���c3�]�b��]�5\'0���ۦ3�C.CS�k�[Ҋ(>{O�&1t�/��ȹ��f�{5'���Ϛ&h&���o�^[,.g�t4���?�cbm�P�%����X��'��ۧ�)z��
��7^��?�{�S?w�)LК�;Q:�3�z:,�13،J�toI�J���{7&1Y?���=�����%1�ޡ���V�p��Vè��M@����8��_����A�V�F)�ĸ�ު^�WՑ���*�.ܙ��h��c��|���DlJ�S}Π��ӊ����?m��,���T�&�%����������{�N�m���#_@Gc�ΙA%x�����6ɸ2���
�e�;���,��u�2庫���������~a�/x�IMyHvVb9�6�^��̨(\��O|�*���t'�l��U���=Y��?��P8g����^i?�o�Xy��3�"aZƟ;XGT-Z}����wy�f�o�侓-��Mq��lL0�R6d	�_�V��1$���i�c�OB�0a��� @b���2 ���i~*1���/�/I�M{�����O��_�y<?�xJ-DP�����qrb�G�ǂ�������:0��D6�:($�#���%X=�il	q��%���}U=�MG*/�~?�.�WQ���^w=��,��$*(?���.�����!Dq�*��NI�<��]�ǥ�T�8�7,F�i�����\�W��x^���+7{&����<�`��;@#��Ϯ�,h�/�s���K@��e���I�6U]E-�pj��a�58^$[-�3��.��e�$�������!ѫ�l�hO��91[=պ���\l�&@�u�2� %?�DX�s���bYow�����H��i��l�">V����B
�+0�[�GAKI8	�m�[�@�Q�̈́�X:Z�X#�O|B�@X�^���xwh��!M���E�q�QAsJo�e/гInv�{�������a�(Wi�5�>ig����}M:��=��b���W>�����Є�De����+TǇ�	t>;6�y��l9�F��v�6�������W$J^7K�W���`!r�Q}��%��ƶA�� �q[���� �A���M)�]�j�v���C�ڂ����ې�oS���bg7���C��|�خJ��}�h�=u?�.�E����Sr��T�ݸ*{�ݿ�%<:j�ܹ�o1i�y~5�Uq�d�D��kf���_�rAc�����śᅟT���I�}�a&|0e����?�6WN�t_Flr����1�y���?��(��f6�����7�[l�Gr#
��I+7� �Vk2~����L)��z�EG���x��W�Ӡ�~l ?�-ؕ(����Η����2"�2���ԩ��a�������(�Q�ffe�A1,�f��yj�a���5F�j=���^�ŃS�_����{|��ҎOj/ ���=�p�6�4ͫ�B�+ͬ�`��[q�MR�Z���S��gt}u�|X��2šT�W���#>� I�C�v�-�r��l'O��__q6V���N����Gw��1��x�����y���pP�Ӝ�鞐��ogiVģ�A`ZڻJ7�8��z^���H`�L74|������6E�P���GJ>DJ/\~6�]M|]`2P���q8T���lF}>�g�����6ZlFe��M�2�´�뿁�g��c�����Tڽ�z^�������s,�����|2��/
 >0�����mp��D��V���#4������ G��4�	�iC��Ԓ��tR�L������P�"�
S���ڷ�ڕ�&��<'�����{�c���t��ð.���Y2C��+r%̇�f�<�0/c����k����և���� E/-F&Pɫ�{:G�ifm�T]/����$_#��s�lBi�[��^���R�Eb$ZiF�(�#�TD�4x��F*�$�����p}��R��k�X���n��E�Gs�w҆�<���=��͚��;����e}Z���#̾�!4���)���	p<�v�0K&��\�M"G]Z���gf��?����%���7`h��.�P����m�ҵ�}v~���B�4�����Wg5���g��|6<�f_�=�i�;Ё�t`W8`}�� ����Y�۝���^f xsL�=��Y:��W�/�2햌nr�r�w���R�A�[���T�b6N�m�X>�6�.}|q�Εf��MPl�O�+�Y���R�oQ�l�U�.�H�����!8�'Fͼ"�EC����)@K֓��lY���q��H���;�^�r?+��/<տ	>Oěb ���i`�n @����`�!X�~�AFepB�04<7H���Fh�ܼ�iC���$�o��0*B`��oScU�<�K�*��8�B��Gi��'{�"��ί�+&B���V�`�j�����& Ͻi��*+�|���4e9��4a|�����������93D��;s�*-9Uܳ���$P�O�����*ίv���!��?V-:Dq�y�0�O�G�<@_>�nyo�X��D`;\L�9����xQۂ}�;T~��V@�(��4�ܰk�>��T)��1��?8kMi��Z8?A����y�D�!8�M푕�4����s�2��29�3L{>��q��3}z����8�-��L�Y=��@>�d�Eq=�BZA\\�s�;2�Zqbc�\�N�^ՃC�.�r�X��&\��ό��Q��@Eg�����DW���+!$1��P�O��9��ʟ���	����q7yi�u"���53Сz�����bs��U�:�sb,���˘\��W����!�{?5��c���Sc��y�:[>��4��Jg)�l��
�M�r���(�����&��b�@2�33�͠Q�Y���!��U����e/�\3@z[�5��4�+��MUnw/>��J�\IY�׃��z6E9<�F}ŭ���2K
��?
_��������#�lfE� #�k�^�7�&u�-�A�{5�{�ߞ�**��rI�$;=;�V�,��Z� F��/Pd@��<��6T����w��p� ���=���)�h�����'�3ٴNr�d��8=}�����Ue����?����k��t������G~�@�`;}a��){พ2ki.�R|[-,z�0�V���ex��/�2{��.D`�6��t�G�.��?ו����&$$�(2���M��l���O��2%<y~�,�s�I�i��;:d쫮C���[(�O9��KW����@�Ԛ�ݫy3nd\`��@�!V��>�XT~p�uá}sam���!*��F�� �B��2.���l��,��ȋ ��§[�7�~�YD���yj��Xn��Q��Z��ct
U׈��.�^S�g?/E����}%�	F��z������z�:���8�A7�Wg��2ݗ�E������d1z���T��(e4�#���\��a��쬧�<�~�Rٞ0e;6>�cO�8	����f ��:�y5X�R9��[ۜ?�%P�}�/�ҋ�	�Ve��]�t��!Xգ�[c�����k���!�th��c\m��	�EE�f��v��2G�R���5�1�π�vR
KJV�&2115K�T]Ϭ#I�������O��PRel1�&�On��N@c�ZcI�)���J�6��e���)��l��"�H�T�Q�V6�`ɼ&����A#��e6�!���<����Q�&;g��X��X�P*�+��˳"FOX�+��b�!L���Րd����(������p�G�.3�Uƌ�0T#f�/v�9�թ��0��|�����^+
���ud�]�,�)z�BOG���^��%y�=��'����i��u߅�*�:���1�i�ŝ�J�Tń����6 D���@�Y����&����+��(������� ����3�������L��DO�%+�½d�W�}R3;c�=2V�|��[���
�c�.�yf�B�BK-�X�А�s��s�+����MF��P����!NK�B������x�T�aӠ�Zbsݞ��:��e�%�;4�p_�v�0��ÍH�X�U���{�pa�jbi#_��	RԩybN����N�H�߼�y���"2��V���ui_�����k�X�]j8��w������F��~j{і����5��Ԅylze�S�{�P�P�9q��x�ۦ��Ɉ��ᶉ�ځhP����8\���j3g�K�c.G��h3�*W�a-W�&˦��/a-�Ȃqm~��CBZ��f�k�⦩E�5�A��10��h��&��!S��q|���t:5Lh�<8���P!�vxӻ��U]{�y�7����ЩyI��k+�&u��o�f݀��,���41�����;U����˴)9�q�1g���?��R��8a1C]����^?a�˶�� 6����WMDA؂�֟Ɲ�-�E"�W������������Ǿ�8�:��=���i�o���������|ʩ��'��,�vz�`s�(�J|lG)��џ�|u\�S��2����l������r���#.[�m9�<��%&(f���]�"#<R��o��X��1�ϥ8}�_'Mf�7��G�M�ƌ��j����*s�PR"3��	r��S��m���X����7��+���3SbV�	{ ��+
�fN��v���/�����/ΐ��Wl����SOP��_��|�)�ف���+t ��'m;�W����Ԕ'[Z���ο��h������)g�,Or�}}����~�]D?��+�fu�'���R������t���lን���< P��k"��i����jND�����$8oњ��ǐ��a��{r���r=�r�!��N���� ��Z��=�'�	��7À�x��vs&u,�Ѓ@��w����VʀS���N�)���V�h��d�C"�ĭ���m����y�7�@�N;��G����(�P�*Ćh�L��6�������;$����ʢ$�;�K�2g~�D�\�qUu�p|�*Q�]�5��8�	D����o�Yf?=gD_S�o�	΋ꮇؘ���O3&2Vi(��:+u$3��&�ځi������h���"vA'�}~,���sݏ�3�!��0����l���Eٌ����]&�9Xq�$f�]���h9`rM3�1��l6Ĉ� Pʔy����(PW[ n����u���m:6;f�q���7�0 ���B���F#�e_L#-����414.�sZ���0֙�`������VWd����kc��N�vӜ�x���
���z{Ðn�R�ya�qE%��r��q�}�,���L�j�"W<(�U��~�]�giդ4*�Wo<k�~��E+NР�g�>b�f,O������c� <�X���� į[�ѭ���1#~	ڞC��x&����{�M��	
&�d�|%�@'���^̞���"�!�|5 �	����V��y�z<�(kN�jj��p��>��`\ g�r��%�A ���y+nM�F���|.���{�I�L�-S�l�%z2a�d�f<��ǋ�<�QxY�	�%�'dn�K�-�P����֏j3�q�g�2ܿ��Y���1ط�Ƈ����#��ʻ���C:f�+ڶ�5+��C�H�ge��������}Vai���j�@ݤ�|Aw�q��K��Ҝ54&�ɣ�����)N5������{����4m�g��(`X�~r�H�H�\�����S��+P�4��ЉhM@��N�*&��o`��L�YB�����b���M5���"��׶�Ҝ��":�� u�'��[U`�_^��>_f�U���\�,V��������}Yu[
�g����a[?7��n������n�r#������F��ϣٮ[D-�O4�'j����9�^�E�O���:mwHeKB:�J�']#��e�	-yGK���I���yg�dm�9z�K'�x�����,<�t����1G�؆OE����2�:�Tj"99bDE�w������m�f��m˳���_m��1�1��Z���G<�@{kK�
.Ԩ�Eۼw�d�ctɾ��%pƃ�b�~Y�WTk��-c��
ED󰘆ou�2��]צ#*�QVK0����b-��*I1Ê	�r�+�i��1M�
9rU�hL8;�;٫�����c�^��ȴ��������a���(�}�FEiAE��h�3k�����faF���M7��Y����|�,B���)>�^�E�sU0�1_�	qrݴC�!�o��Z�2�%GRs]5/�X�]F�&>�����AX�M���g��P����[��:?3YLt���:vH{��R �C�b=%VQ��sa�^X�<U!��a�o�c������9��3��6w8v�"�Q(�\�B*�V6�\y:�ߗ�#M�o��4�>���ګ> �څf��� �����k��^����MW���p�N߸��n����A��Z#����8���ԨbFFn��mR�y�W�ǵGA� �}`���N�q�R*���L'5U,�ċW�L�ZiM��wծ#N�|���f��*�j8���ru���g�����ɚ��T>n�\��;u����q	��Ǆ[���_0FZm0��K���	���:EH�Y�G@�O����]=_���T���m�r2Z(zz�(E����>��ִ�o쨈�U�*���B ��[�lk��r4�-?��t��8�o��+'z�C_<�3�� ~@t����eveP��Ui؊#�;��B몀�^�-��Y7�:~<_G�E�*+�j4�G������s�~}r5�A� sq��z�������[��I�c�!�vhJ�����R�B�4��@G�c"�f.l�����jUbA��ݱM�����hz��ǧz�t�E��醧�N8p�!���ud��s4*�}"��b�Y<�6�S��`�����$C�(�JV�#�QD��e�TG=���W}P��tڼ�����&q���u��>�&��ڞ��dY+�|�)����&�D�_�4�L�Ԇ��9{��k��'D�	+ۼ��4����0�~��hd�u���g�{����xD�w���`j���0�(��~�޴y�Cˡ�ތ�#�w8B��!q�>X,ލ�Vz��������O�V�P���v����5�x�ٔo�rY ��&%d��X�qm/4#�PԤ[�����������K�~�V���a ��%��f��f�l�y���g��Σ��TR�gE�.�m��-�)���M�u�w��Ix�+�*��l�+�iSD>{=f�X�
/f���V����#���Ql�>���6��j0��5h��E�~��a�����z�W�����M�f{ݪ�JL�tqp+wK��]��觰�:m����2p�H1�q!s�3!9�����u�y�k�/��XZ,s_���|��Jʋ�k]5!�8�`�e�Ì����b:��~'��Nu����ʍ�ڻ�(D�
�8�x��܏�G����U��J�Fa	4j�i�`����1�L�f�P�Z�YOxĘ�B'�?���,��S�D2HR-�_���0�����a�F����jn;�r��~ʊ�Y?�Pފ��#�J�&����pe�� I8oo4MkRp�;�4��,��S���ͪ���l�����Ѭ\ ���Tc�H̦9+�R'շ7�����8���Ź��A����A�2(���F�\�;��!�4��ܯ�܋q�O�%VR�i&��!1D���~+��z�9���i���j9��_����V��0K�<�3[�9[����� L0���q�r(ڷ�m<t�φ5�=�!P��(gN�^*F����d�GN6ĺ演�Q����w˧�ޏ�j�Ӷ�Q���4�ph�L ��	��w��1����ݝ��"��.Y���$UL�R����O6߸@�=����X�˖F��@���R�!u��v�+� ��x2���(���g�͸ �qZ��P��8�	ru���-�#���~�#>��3�jC&2�@ӟGv�C��lV�w>����5UM,��+�4�M�`�h��R���4���..�I0f�?�,nT�ϖ�>4�[�<x?��}G�%U���0�D��0=馒����Y�4��t�lF������ ��k2R�Ԥ�^����GV�~���O�'�Ŗȁ{`������?=4�RzخAI����\ZCEj�ϔKϡ���_�sUX�$=�]�>;nfQoP���({��܀�l�H��՛�w���o�&��_�Aq�[�н�Iݟ��kxG����wi����F�B��KIh�o�S�Fo�����q�7xz[r�{k�˻N���@wN˂�+{q���Oui&��*ٸt#�LpŬ/���L�5���W��xبN;�W�n�'��*̗���֞�����1�*�ZnUt�h�ZӰ/ǳ
��/R� ������P$Ɋ���d�f��,K��Hj��Ll�rQp��:69������gi�c/̷�Z��K4*S�uוp	�땮qY�}kϛ���:���dD	l@g���#��E�fq��Tύq�s����KU'(���Q$��t�zws�"oh׉��F(V�MC��x��j����+Ȗ���5�j����?s����hu�,�0���=��\}=��d�
�c)>�&�����d�칤�]mҐxc^��V/tE��}t���aT�gn��~���kͪ��`����X����h��|��QGb�{9����E���cE�Z=�U�����Ø�C�C�e���K���k�0"6�d�}hʱ�}��5u��TǕ��G��\��A��K]��=��h�]�l�E�[_1+��Re�Z�ݢ�]ã�m=�]�,���
��]|l�coyiJl��	ǖ�1�VN+E����;�7$��٣#�&��`J�!bh�^���`�����IlW�0���W�3�ƺ/��q�b햢��ũ:<�MS�I��os���L����qFv��~���aDmlp:�Sۊ�pU�0���U���W�NC�d�t>I,�ě�����j��usi�O3a�1�j��gc�Z�Y�y�9c�U��mh�!�7 R�e��v��W*��<���滻J��\FrR���b/U�����*d]g��M�B(�K���L������s��'�(�A��&��=�����G��_ys���S��rW5�]+���e�J>��vI��.��MJ͒JM���F*R���[���f��+d,|Qee�B/��=kx�]���`Ѫ���9��uCX߅��k1���-y~�%k}�=�@�x�!p9�g��=��́���!��`�����'瓮�_�x^�o��@��'ұ;�u�D�oxS�rY�k�0%�g�^��>�h��=�#.U��_ay4�}��R��F?�J���}��rq�D3�BN�:���[��$���o�E�����&��d ���s�z.�7,"��������Ie�9��J2�fqLR��ņ�&�:�E��{���3ב�*���ĭJC/]��fd;��,J���\���
�5����{O�H�%>�O5���ҁA+�m�mB�8$�4�e�*}�j+�)����{��s����g�y���7��r=�z�S���pl�rϭy�z�#�׻F���[/�/f���R��m9[s-&�1��/R�%��l9�D���%
h��e۰#�u�kB��t�reM}[x5)q� '���sGӵo��R�n�|��"��)�{��;$Ӷq�m�c�Y_A���F������k��v���O�nxLg�m����"�3�*1�Z a:���I{�L��Y���kX�5���-�b	�	܃44�R�<R�׻�4؞�G_������#��͉�a�;̘���l4�ݩs$��kͮɾ�o\��� KR����v��3T8D�m꫏�Akc��TE�n�u�}�@Y?��}�� y��Z�4��c�)MG�ї:���=\�c��J��eV�� Q�	r�뢞��UʥOs��꿼���.Еo���z����t&���9/G!GJE���$�cfb�t㻗��b�(���Nɧ{�L�²��$ط2\{��	X���<�8��C��1 ����J Q�L7u�_�n�3 d���C���ݻ6�:��:���0����<�K�x9��7����w�jZTn��&�9踰a��0����ǋ�T1�����@|���8ːy�[M�Y����g:V8ݿ�f��F��[��r[�G���p��軨�y��˷����QP�ˆ���mu�3&Bf���o��d���0\A�΄V�@Ƨ�����Ӓ̋>Hg(h���Xg2�ix���}DO�4m�x%�̌H�����]-�?�Idր:NPTP�\����5�l��ѠC�YC�?:����~ޠ����u��y�y�8�$�;�+D�8����c�a�(I�h�c�;��r(Gcs@�ĵ]�+���%�`�'�>�#��4ٮ��G=��h�W��Ψ���~�~kW$	�q��x��.��� �m
Q;�V4}��,Ű�;��j�*�*��K�I�����������?�X<s��(�v����ʻ�sBA|���1��oY��}�'m۷2��f�V7�43��X�m������R��y�{�tbh>�CG/DvP�C�M#��O�at��dy�N<�ȋ� "}���L}�0�)f�� ),��0:��6C�Ҵ�N�!i����Q���d-�ؒ��x&~..]R-��/��e.����b�[�E&+�{;۾s?	I7���#P�ߡp��'�{��;�~,`x������6&Vpg�F�����\Ы|f��3W��؀��n�il��Aư��b� �j���f��k��92F��.v���ya�#I�g��m��_�*�����P�ߕ��a�^<�89"�A~*��J_��bf�Qҧ)[�i�V�+3*�z��*O���2�r��y��m�i�<,��%�྿7�Po�`�1(��O-S/�X��v{�M�]sC�zw5���Yt+7*Hb�㾤2�À�O~ZЃ����m�>%/�ZyZTw)k������K������j6��~�~>��b�@'��35��hGAB���ß�r�k� ����N�h_D�~m�g�"�$\��\�/�A�I=���\Da+���������Z�W��%�ʕ^:�I9����ȷ3eE��6�lRҹH�@16�L$�P��Gn�?�W���kh2A�^�g��$x^7!�&�������� B�LjA<��"R{^y�<��<N�U2�z�Ê����ɚ[���V�~:+��}|w�1���_ݻlߜ�XY�B�#A�,�1���'?�I4�S֝��3#���}�ヶ��k��ֹ�E! �T��?Th�'�/b�]�����R�*Vx��T��uXB0o~ ¦q�"5M�ɫ��os������%�(�Y����FU�����/��y�r��DѢ�J~ �t�{=�^��$�	��#�_�� ��E�ơ7����ҽ��#�EFn�ɸ	z:RU�oxx��X�?�06�oZ,4p��XY��~���	
�Ӈy9�%HkĄϑk�O���79� ������eK	��!Reo��a�'[l�]"��%��$�(�)A:�%����9qRl�{l^,��<r�-_v%�R3�J��2�╌'U�Oבb[�G���8�
���7+�fء68�ɅĠ#)�B��2L�6e�R��}�>Q��"�V��g1G�3I0f߶�qݱ�Cς�c�7VOS���ŬM����cy��Y����!B���ɀ�1�1�����v�����ro�Tۧ�����\�4�Ut���֣�g?��?�����\#�>�9� {���K?����s�A�����`�r��u��� h8U���)n�Y�N����R�]h�*��*�L�+�m}5���+�_��%��*u���E��9F���y��a����L.z�Yu|2fͮ�A��&D4�Z#�)�<"��䌦����'�&�A��xX����oӑ���I�FB���������5��|��0zw	t��7�N�m�{�仐Z0Z���h_����;��w��`�G��T8�O��������rZ����c"i!X�����Du~�he|�T��d�E�3\������eۏ�K⫻i�g_���ޅ|�c���mqY���Ѵ�>�*8�qX�ȠZ�f�|*Ԁ����O1��Э��O&��qᅬ!�^f8 �b���]����00�xՈz&S�HmXkU��~���w0>%qP�U8Q�.��[�*<ބN�v�Y0���xdg�����4��#L�kh��.�4����#^=Q��6�
9 ��o��L,�ߙ	k[ͳ�Z���l�CIK��]��=�zN�V3L��<# �6����/}!�(�QN�R�Gj�4ǟ��n@��w2��
�,cջM� �cRxB�ݫ�,R#)��W�m�����}bu��s��(V���?	r̴%�=�1�n�&6K�_��ˆ�=�6��Q� ��0�����%XĒ`0!W�b����[��G�Ə��=�5=&��
���pL��}��a/���!�b���H���/(�('�,d<��hϏ8�0�b�2�ڶ&dݧޛ�s@T�H+�$,t��2K��G�X�^EMcFv��d&2ۂ�eYM�8ZI7=In�D���7,�'\KXŐ��qa�6�^���V���.s�Z���t˜S}�����@��#�b ߖ���it?�ca�cp�_�D��"Q0�Ӏ�*�DE˴���qA g��@��a��Z��Jd`�d�X
����bP�W�4�����2�!H������c(��hS��+Z3q�U����� w@��n����\OY�LADٔ[��fQ �L�Q���OU�2->�ӅvvW����4�T�X�Ey�۵�F�  �Z�v��V^���Y{����Wsº�����
��xd~CP����_��o��%�y�J��E���s��t�Iv�'z͍���f7����,A,��/���Dd(�AA��Z߂~�<&�D�%5��<��|&a�����`��]۠�2޲�y�t~j<�9~��G�?��!�9�Aa����@(�L	�~���g��:7L�/�����u
<
R���
$x3���y��Vt22���KVy}j���-[��p�p�1�Ⱥ�{X��֮;2��<�kj�nU��=�=ϩ]�O�m`�f[�n�]#��Eg��������wXc*�����!������#E���	���z�B�&�C`-!gT<R1 ��5��>���;�$�9x�+^a�������L�=�8�ą�llv���\�M��#�o��j]�!2�r��R�����G�M��N�`3#��f��M���|��ށ怍MYo}�rJ(�E� �α��T3L8��K_�R�`�6�5���aY�z���\*[<o5ptʔ�n8,�V<�%���_�<��4��7�:�vf����>�-�3r� �+{��m��͙�O���3[�G�-�G��jj���P���d{hƼ�E�r�adF8�9�}���۷��-74y_���}�Z�t{_Z�u�Mo�2	��]`�Lf���X��h�Vv�5��cc��z��|�� Z���B�O1AM��!�������P��[�/n��-�#��=�	N�t��!�ʱXt�1���!!�b�ϳ��*��k-Oc�m@$��!$��eW �to���ޏv��ɺs��/��pZoI�4�lr|4}w�W����񬍏��/����DBXR��{3�\����,��莴Ӈ�w�Y}")��	� ���Ζ'��{��~�j�P'��C��/��,Yk|���kr���it$��);�3=�り��[�¿��7��u:N��{���`/������$O��g�����=��cNGcA���:�l��5���Kq��|��ڱ���Vڐ�)�zc��}��!��s
�}AG��-��`�}�L���y>b��#.�����0"�0B.������9��KC��]��{P��W�rn?�!��7�e�gX'S�j�6h͵����*�{+c�����~���dm*��]����G��~��Ie̜Y���=z\���G��O"�/��iC1�\��U�����{p�~Z�>zZ�s戮�?fc�۝�99Ѱ�;��W������^ ���[y�,S�L�{���66���$ͫ��t/ɣL
��(�t\#��N^��K�FQ��=���	.���l'	��K;(6����l�F�;�jW�ȚfRV�&�~����g0�>�\;㌳|--_���~�/�Z��[=�����z�pݢ���Kie������<+=��/�'�x��=i�֘�x��~���i�G���k��u{�K/�3�8�'��LJ0^%6q�#�8>�h��y��z �\&kQ��9F���0�s�(x/�|��f�tfs�����+�'E�8�<		љD�0d��#�,�ى���Dƙ���	2}�����"h.�c]����'�*g�9����SXO\O�qRP�!�JO��ݺ�lw$���k֬����:A�48ɡL�v�u_K�`�v��Q+�j�Z�CIy�%,�q�fV�U�
��u�s��DY!���R�>b~���M�/��j�aOm|����$�������Z��{vϝ��ӛ��W��5�`�,�+���6=����;�\�4�^�[�'ּ"�g�y��Y��v��e�n�d�c�����Aa��Z���i�sɲ۽{�v<7f�z�o��N;ͅ<�:mv�8)��đ�O�=c��G}����SP��^h��bzc��a(��"E6&�D�+:^��oi^��
�J(K��<���{��X4�!�ň��D4}�<���P�U����,&������,�邔�o��	�$^5���=��g���V�В�[�K�,K�g��O�ã�+	҉�,ڪ������d�����7����[*��wK�Sʼ�bm{�(��L#sK�Z#����#���_�`4�~ޒ����lI�'á���NL5l|l�x����/��b�y�a�=>əg���9`�����F=��Sltt��4��v;��c�ϱIP?bc��aU|a�	�vW���^���y�l�&y�{��]�轉r �o��o�k�q%��_~���D)�S�_����z�������S �K�ySB�	�L�
D^�ޏ�:#�^�}��)&��K�Y��)DhH�9����~
$G��5�ZP����5�,}��r����j(�e�A���-]���E�7�9� `hi��p�+4iY�4���\�w��6>9���@s�.���|{����o[���M�Y�E�N�sK'.�c�ȹ^}�7/c��/��7��G{ ]�|�z{����y1��Fmْ��s�6Wp?���SN����8RJ���;��x��"��^��zp	E��&�k����㫛6=n'��Q�  Iԝ?6e��
o��+��	�V� ��!������+^��g�@�cA��Dt��3ͭd��1��s��`},IA�����;���nd53g��&�R�c<� :�,���{#<����^S���XF� ��^��cnH���J�f�zbI���z����FV§�,ٵI�Z�ɾ2'Tp�����xF�M{?aɲ�~��oM�=̓�H��MP4��BL��t�������[�P\�Z����˿��EO)O��}��=��ԭ�uĞ���C���ڱǮ��kץgٲ�RSHG��/������?��O�|9�c�Gy��]s�=����L{K�]�¿Y��I��o��>�����b=�١���1�oƴq�&���O�p�|�^m^�
����GP\w�u�pp�	��A��c�wdg7�e���)��i�,Y�9FPJ����`+�+�N�U�Gʇ��U%�c^�6wL ����v�9��>�����=|c��{��v�c>�l���";e�J���,�Z���w��$�̂�N.�'y%����+��!��'��K���=�c�-s��R�J�����h�t\XK�����+�}��;�<��_�U���߁��xd�>�{�;����Xc�'Ň	�Ï�pX:��k}�<���#�<˕����ֻ��kiM4m��U��bMD�g�߳k�E/�{�RK��N�/��/fN�&βɫU��M��L<15Tw#�*���~�!*7��]�C?��ُ������U�)������o~�uW6�V|x	��M�yC�K(F�����G e�g�}U��0�!�!(F8�KxpN>ˉs����j� ��x&h15��"ry-}R|�+X�E]P��-���پ!�)}���\��,K�VYe`iV��<@\*W���=͖F��e{���k���L^t0��̋�5�I���l`pvڵM��Gg<%2�.��b�l��̅�#HX��G�I[X�R�j�����x.�:�H�7�CN�����d-M�-}O�^�ٞeH�B�]�¿ԍ��*����X�: ����g7�p'����崨�_ZN�C�)�Sw�Kբ��Ұ�y�L=�gV��63������{��`�j�� ��m���C�6�K6Y���ñ��?��O��uϐU-Z]�dp�^�7��ω�zXj��y�!�����*՟s�z,�qy��g	l��ܛ�N�.���k�\�"8�S2��jȒ�a�wZ}����R^A���t:o١���cɫ~����d�[�:hO<��Tyi�HR,��Z�]���\�YO$܋�U��F�9w{�x���퓶eێ,�ײd��h�;7Hs)��%�!N<�g�<���c����ەQ���	JY���+�{/�rqT�Ȓe��z��}�6[�r�mٱ����X��?MvO�<�Mأ�<��Q�O�Y}hZ��41#Vo���I�Q�vȊ[�{ܶl��欳�*�Rzy*�Y,,=6���h�(h�U��%�����C�YA�K/����R�S~A�?C�y��emɲV�%����0�����<G)��ȸ��T4N�:k
1���m�g!l����E0Od�Ha�}����׾6S@�v{S���ط��9$3U���-��cTbw����{�/�R��ozf��6����$,���t/O��q��$�К�q����K�+��4�7���j'�u*���i%H�^�mS3�k_��~����!��!�0(š����S	���^����d��x\�5�j������������gmbr�ο�,[vH2PmԞ���m����M�:)�4�?����W�>�,b��|�N8~��%����`��w�m~v�'bd1�J	����$�e�~�!�iXlR�{UeѼ���׼�5E/-"ea�qם�����w�/���b���nk�^�\�1cFA�Nn~dIȃY�A�J��>:���]*��f�!Ų!�.�Z�*8'�qxZS|E �q~��
���.���u��攋��4#�gF�TBV�ٰFS �j*F�ߔ���>�{d���`�Y�9��\��_~V�� u�/��H��V 1�+��d�`(�����v�/���7���������=H&�u�]^:f�-v���m�s������� O�֬]jûFl鲕����;�زQ{�)'y�J�����{�"ٞ�w�V�|`
���/�������ڹ��V�X�A��?�v�x��ȳ��5�竖���O{�����t����n!)���f�����G�f�����ۋE<:8vHX��M�9<2���Z�I��Z����I�߼�< ,��2�ʊ%H1��t}X���Y7���i���~,�s�<M���m
�CP�9�
�P6 K���R!���� �(2V�q��hgҔ؞`��d�QnA0L��GP6��J���������B��[@!R:3ɽr� �m\ż�H���Y��{��
 ���y��fB��Տ��Gp�q��e�t�HoH�߿�6=�ɦ&F��Y5�Om�dK�bkWeW\v^:~m�%{��-�u�D��c��V���0�)�΃�~�;��;���68�o�#%;��b��m�=�̟&�1�S;����/��ի�M07�ζ�~���{��%�\�A ��x�^np�7���H��3�����CPV0�1�X*���rW�f;�uZ���`I#�# �sqNA>���'��Pք���
^T^�M�`
�F�c|�-�׃����HB�\^zd�]�Cu��$�"b4��HT5U��,����e��T:�j�2ku�Y�	b��
���\��_��@��h͕ 17����+#����}
멼6�!�Q̳�#5d�w��;~�*k��ǜh��%v����Ș=��öb�!�b�Jמ�^t�u�zOv���w�{]R��ҵ``�|X��?���ߦ�\���j؏�3_�o|��m�в���^}�v�k^�Y�XC�w+gk�0, ������X�:��l@(�#��f0-66�~i�}pt�hl`6�\|��W�R�� ���H��Њx�b%|q.� C���C�V�`����Q�]���cbd��^QQ1B���׃�y{H1Q�2��}��z�R�S
��5������x��&-�
�ߖ��
�>]h7m�׳�Sn��f��?�{�
Q��r� �4�����9�������x�}~��󁒅�)
hdW)��*����y���=j+Vn������7$I']���G���F���/����v�=^�F��}�.~��*���MF�ʕ�=SʉA�����ܶ���.��O~I�*��<0�ԅ���pM�5��޻��	"�N�j2�l(�?�я��� Y���{.��U�����V7�F��o}�L��_�Ln�R0@��ɳֹ�{�O��;b���� ,tq��W�0G(`�5BT� %֮����`ۇ�r�b&�cP\��(^��W�ҹ�%%a�V?�60���<R�5@���D����Kmf0�C@y=�v\K���;�tx)�������f}�|�H�-r �=���Tn�09<(]�9�F~^$L);/�9^��o;���]l�Y�k�C������u#6�d��عծ��Z��G7gl�ь-V��3�X�¿�h:elddgf���&�s��o?��v{��G�\
�أ�v�N�e$�fvo��6{���{,�F�SD�����?�C��h������KH0x������_��p�YXjxp,�P�U��SO=5#t����'�E#�폘?CBRyZ��Ǆ)�}h�cP] �t>����G���,�I�F�JHIgA������>Q,JTV��;:��l�{�<���e ;���ؙ?�Y��Z���]�ᡒ��l��{��b|y�f?.|N�X�>�6bM$����I�p>���"���gV�����x��<w��7��	���o�=���u��?~��vc�ݲ�5��!�n����o۾��ȕ(��G���4�����7�X�¿U�N�ECg���W+W������2͎����h��@ڠ�b�U�z@ic0�X]*��q��;������)AE`"(������2 8�`a������M&�Q���+P+H�y��3��$P	�ך`�F0 x���q|��W0v�S+�22��Jb�7V������J̍TO�Ž3��4�P�PD=�{�k��_�F���t�l<��P*,��&� �C� g��A��R#h9{�����,���m�pD~�1��1xy��{���+	�������A����	ni�3��k_��?+�Eo՘nb��ݶcǮ�HH߅g�{x��T�̳Ƣ��GZ�Su���H��#ɵ���0=�:����i4������d�Q.��=���ܥF��D��44�����C��O��Ii0�0��#���M��N�'V��KL@��|�`�`�tB[X�k�軕���=�ǜ	A&*��?����x\k�vQ/���:��(�I�3ޟ(��B&+�*�C,��;dH �r�:����J9w
�%�Z>
�b����l���P�]�>?��`l���<���i6
%��(XS�\�6��9y/���l�|9+�9W2W��Ox6q9�}��H�s�4ʘ+Z"��K1���z`�(N
7�����=�����q��栘�A���G����"T��0XC��Qʆ�c+}e9S=�S��J��l�����d�Q|�+��E���z��ڸ����"b��lŅ"�7�\��K�D���E����BK�Pcq2Q�|sV�s:�>�wxE
^
�%h�������l��#��m(kz	d+�h���E�b09���e�k>�<�%)��ȥ㣱 ����ܷ�T�,�u�NA���	���me4�y_��tEPˍ�z1z���3V#.�>/�@7�̸�*<s*�:-�ޚv]{;b�yUڧĀ����@�����1��`��=�{�̣R����{��E/�{|go=���:Ӛ��6��?�y���aU��� �������>p�c[m4-�H-�9��mp�Z��d��ǾЖ�(��k�z�k#d�=�Ȣ�A���	�U�G-9x�U�E�by���Cשu��v�ɳ�x�X-�	%Pe���B��!ڦbU�������*��"�\D�z2��s9�`�}�&���aȋ�E�m�Iq�kjgHO�=���sYM����ڰg)�c�՜^uS�o��ٵ�bn�*Y���y���g3��s���]3g�*F�gV���_��{4g��sE�\Q��C@������r6�,G~�{�.J^l�.�@�p�v��mp>��N(`(��B`b�r���c"�Y�);ݫ��7�����b��u������0�O|�^�G���m.���:�_��`4����r�3zF������3|�*��8A8�Y�4AN�֕
�EA$�&!��w�N~9,�}ҋ�O<+hܫ��")
	J�U�b�n�2%1��IyZ���htXx����{�}�D͌*]��_aD�b��wQ?�)�U`����^������(�p�	�qi�,��YQ��ͭ@��T6%���*�Å`.�bC��Ҩ'X����õ��׮T�,��χ�/Z�P���8��hY*Q}%��g(�B0	�/���S���΋*M�0�CL��9kPP�2�uY������Py�����0�C�`�x�:��T`�)I{gEC��P�Vre�r$�cs)<�K���>JvblԿ��#��ƾ�[�x��5��PW�\�}�'�۾랻3je���3��"�.���yD�;����l��!o�y���G/�f�8��6�bD���m�շSC�J�Q�`�K	6Zp��TS�H6�m����h������X��}uǠ����Z����9����{#���|
�	�ݟ�{�C�A@$zqR"�^),	�s�~�o5fU�k@h��#HBВbGz�N��ۇ���w_	y1�$�4���nCumtm�l��~V�.�1R#���l�[]���%̹�Q���L+y�*q+�F2���^�c����X�¿���L?�g�5�.�Y��̔�� WPM�{��e9�/�_~Yb����f=��n�%��X�,/p�a�~-��u���L��r�|׎�UU�.s��9O�%Bϟ �,8��g�u�c�	�^��ye5*CT8�����$o	+��V6��:�X&b�ț��8ߍU�^��"�7]�O�S�A��P�N���X�VJ���,"�:���n�R�i/��k428�k5g�Y�	���3�� �C����V��a|1�C���ǿ�س��L	�1��o�/{�m[3=���L��5���Fĕf�`�j�ֺ,5Yڰlq�%P}��zo�XbX�.��r�^
v�M�0�F�L���k�cD�������� Ās'�R����}|��T�-*{�C�,oi#{GX3��n��_�ñ�,)�5)%� Vf0�ٯ��
Q��x��̫n�W�)�:8/�'�*,~h��>�=�r�6���a���O#�Ә��i�hOkϪ+\�w]�n�gX��sؓs�\ا��nf��T(ɐM�H�|�g`��|�X��h�S��j�K�F�/��P.qt�5�����V[xE����,#]�R� ��\ӔM��H@ĎO�4v��=]C'��=Yt�0�|C|�j�p����eD;��g��֊���1�1� n�Ź8V5���9��5[��,~,v?�FLYE ��T�?*w5v���X�3i���"���nR�P �:c�X������in����U��e�4��_�1�O�gQ.�Oĩ��L��֥�2
}]���u龳}���~n�Cy>�d���6�!��"_ �����@E�^���}(�P�fV�X����f�)�x�q'dV�Ĥ�G�mٚg�V����%�!+�����Z�F
c''��-vX�q�j�+`k�hQw~N���3a�^�NX�ҧ�PbP�G���GB!2g����PB�y��+K�90����a%_͵ܶ�έ��3W醨�Y#@�
��<�	U�Gx2��O��ד>��se�F>�=q�W\qEf�4��`�S������z) )�+�9w�~�扌d 73A��׭�ViZޅ�����K���~R�=8_�z���'��1���^�-҃Y'�p�y��g��@V�i��K�����
`��V�'C�4��7N5	��1�:'/y�K���3���)�:�&��d�y���'K^�	.&.��O>�j��~{��fcSD
!�[����`Y1�Ŭͤ���)dU����GL#Y��F���QK�G&	#*3)C	����!O#&��߅V 
�I�<"�F�Ne�
��^P"�G�\
E]��1>7�^BZ��V�̺&���:G������JT��!��2�״6���:�����9���z
ȫ%�Kq�n�[�Qݓ�Kk�כ-���u�s��j�+�"3$�5�2���G��^��N8�=ϥK�����n_?��Ńv������lyY�9�t>p3|���U�gVOQOG����|�7\��H�HL��f��V��&k��u�i��op��L:�~��~�7��_���\i\{���]Dlu&�Lc�4{�N7d�kX��%������Ɋ��YC����Z�Ŏ����N��ڬ�.��(����u-<�d������,AS���z��u%���6��/(2zCR���o��0^BK]���u�μ�V�iD���T�UDl����Dh'Z�b��we�f���lC��O����~ �uZ��W��(���!&���d`R���3�p�oȕv53��9�l����䦧�_�G7 �U"�P	t_Ǣ�y	�YI!�Ed�j|/��"��񤝫e\�qۼ#�j�e98X�ɴAN9�$[�f�O�����ª�P��K�����|�7ۿ��������^�Sة�	Pa�sI�P	C_MA�� ���1K! ^��C�G�j)���'�
�ٯ�r�3v��,x���_��(���Θ��/
�s�]�ys�L��zI ꘨e`Ȼ�=d#D�s�L*Qu�����y]�	����n/?�ZPRН���Q�1`�ƺ֩F����Y�KAc=��&
\x5Z����4��a��⾋Ɣ<���Ø@���կ����J¨lN��(�8͂$���ڵӖ,�����>�[�/|�Kɀ�ϖ-Yj��#��q_Ǣ������˽�����^��+��9�H���n���Y�W�\�=8O?�,��<X)Z+^�	D)<��#>���_����|�#^��f,���� ?�5��׆CyQ%/C�v(�'�9��~�(9~t/j΢���5����lV,,e��������Q�Œ��$ "�����qi.��z�h�Ȑ0��=�/Z�<�JR�1�'��R*�������R��bs�H�t��Z�E%�EZ�s��'[U+E�YJ^�+���q�6"�罠���@m�7%�̟����c�~�^ӱm<\0��z��ב��нy	���0������R���7�>	~��~��6nz�n�����;}n���=�<[��P'�,Y:h�~���_����^��A��v[�¿Ճ�59Q�`��]#v�1G����d}�U�?�arٶ�q��Yv
��/�ݞ|�q;�e�Y��RW_|�G5jg!bI���p!I����ۇ?�a{����3ZGmj�|�6��(l�}"@X�����k\�h�	o]�g��9Z�q=>��X�jT@�8�\	&Q��[B^TG0N~7z�Xx��6*�X/E����xu�*1���u�־p`�S�]T�A�-���y=Blj���C�3&�˜0W�a���=�X�ū 2ǣ�E!U��FC�q�Z�_/��@�+��(
���e�����'wq-Y���;�1��3'W"(��<m۶=�s�C�����h��=�y�k�A%��g��w���2I {n�3v˭?���m鐕�%{��_�5�����^w���V��UW������vNI��Ƣ����dc��\ȍ��N��m|�Qk�ǒ��O�t�UrL��o�޴�׶l��w��}�ݑ D�M(�#��F�W4<�dY�
|F7�׈L�N�!��M��T�b�Y���М�sa��@8F��x��
�,S�	�X$���*!#Ꟛ���D�I�="^�Z�RFX��	<:���l7�' K[ޒ���.��_�3w�F���������q��3��U0a���jq]��՝{���7�!�-4�5�>��Ϻ��� �8���q��<��Ig������ܙ�+�?�
�zQE�������o�o�q���\��1��?�>�[�y=��Rԭ�1{v�S�s�6[���zkmbr��Z��}�����ˮx��AA�u�v��?rJ�/�K�3&��Y�kIz��^nL$��u߽ގ>v��o8̞����L�?ɽ��)�oO�J��Э?�Ņ��ظ��8{j㦢 ����)�.���B�_����n�tz	8Q��^GFE�5�G�g)XJ��\��,>5���*����BB%$T�����e&�@4Eᘂn�#��`�ApR�k��vX��/4癝3ǡ����i�iw&�u+w���Y�\�փ:o���v*�^�J=(ʔ�����&R�������|�yWp;��el(�4>9QԧaD�c�F��@�ր��+Z���״�bn���]�J��v:xql�O!�F�<CFRr����oذ�~�#u���o*�;��Uo}�-Zb_��W=��o
k�b�z�+���+�mz�qk��؉돰'7>��~��F&_���-�����V;�S�_���Jo��hvx��@�������;��;�V�\�&��I_���u�G���6�`�)X�� [��1�,(K���kXO?���@*��𖷼�q>�,����?m?���E@/�ᴐz�N�Yt�8{W���B� ��,�����o˞��>�@R���^�Ғ��+!
S�uH�I���|�>�];-���k�gAO,�p�^Z�zL�L�Z�+��|�[���gd�Ǻ2���	B�������&6̹+�r�5��	2�ٹƤf*lV.5�&�������A��KVt	k_�����s�X�b)
����?���Z+���~��N㦮����<�����{ϝ��C�@J@�S@E�����T� ƭ�2h��� qd�	':DM< ��g6�A��+Ib��v�����R�d�?��S��-�m�&3�Y�T�R���L��h7�@X
Fbc��	�b�}�;�q� |�w�w��?�)��Ul ыJ7pd��������H�0J���	�$�)��<�J����ıD#J���P��I��@4��D.��1"�U�
���+���������;Q���>fbGVH�̙�ye�:� �ǅ�G9K�k��(
�v>g����g�W+X'*9-�W���fce־_���ݳ�{+�L�]O��:��ÿć~x��n��!��e�ā~YGxyt��|k�����m���y�!i�ҟ���N��O�s��=���o��VK�x]�\Ǣ��L_���0D��rˊ��Ov�����I�*-��!��X�C8��t�y�{�:��ƥ�'-ߨ�N]{�L��@Y�)��ׁ���
03x��4���V=�$P�(�)I	+}w��kr���B�\��b�;RW�rHiʒ�	Uz��+��>���6��ˡ5֔<��{���k� �
d���?� /�Y�����%����,�)gP� a�
���Q.�z9Nީ�J�=�L[6� �`���c��BI,��3�bє�u�O>n�F,@�%�� �D���-PE��O�S��4��i}Y����<:�ÿ������OL+s�)�ۈ����i�>����l��z�ȏ9f��t#�+K"�L���db}9������H�Q�H���l �"�;�3N����Z�!��|���ǚ�lv�HmhY�F��1�����Y��7R�$@�����R�n�SѱN��G^�8�ԘG!J�1����������6S�������P�q�ְU���yMA^�Q�C8��"��d2�R�z�/(���oֺ�ː�I�����?��X�)L)��-TF�c���$���O�q���-�׫^~�S�K��p��ۿ�A�w���M��w�y������>�o�!���[Cs��_s!�m՛S6���Z��rr �ג���2���Ĩ�5�!f��9�E/�ͺ�wgg3`~�a�j�a�;�OѶZ�VV����Ln��'m�ݾ!�p�$&M�*�t~YbJ�<� �"ZR���lC�����`���q 1��6	l,D-N����q�����=���c�^��V]A��y��"�^����%mJ1pH���+Ȅ��f������^�g.�_�M=7��
ݕ��uQ2���Aq��0ψ��=A2~e�j]�X��o8Ya{�F#�k����xĠ�����i�=͵�Ѿ�Rkv�L���mHc��{�s���W�ʧ���8X~�m���<;�XO��������X�3C�������,����lt��ɦ�|��>gcim�Tdh�
�&E2�\�¿٣����l���^y�����s^�lOۮ��l�����F�(��Z�R[����a[w�R��#I�[�8�2�#�KO,�E1(
�ن,���`U�W�_�;���}T���X���r��bPL�t�$KV�
���A��C�Kx�*����v�������n�M*�D�LP������υ�h��f=��1��
��2�A�1j )���`p>QL���QS�L�Ab�b���s����]��cnj��r�v�ry�z��0�-�=�N�n1�00�{���!}�!;�%��3���۞�F�φ��:��4�v�I�أ�lLϻ�pF_2F�3��w�O�&����;��9�i��g.8��$�WZ�@5�W#���:�t�?�g�Ɇsp)�v��.*0m&���l0�?��?م^XP�b���G{���ͯ`�\��%p�0�YE���>��f�9����H��s(���C�0F֢��V\��͓!�\�AyX/�>�5<��"��h���6?���$%X��P�e�� �,ƙ���A����H!w
"�Oтǻ�F��Z;����C���ľ�,��̚��o��33��o�s��&�^�9��3��潔@l���-oՍ��z�a)~�'��7���>��[�;e0�&Ӽ�\u��ܽ+}~�m����J�犲�f�d�Ye�^v�{�z�<{�F�����/�Z����'�BIf�;��~�n��&��5�Nx��:f�/͝���'7�3<n�rՎ8�(;��uv�y'���MǺb�p��^z�M7��"�gS1�K��B8W���Eb)0���lB9&����|�7C��K��{D����uQ�-o"R�Ua�XH1��x��l�wO O-��cEHE�L	��6��Y�M���3R��m	r��P�;��g�a�8����D&�����W1�"~��dp>�����`�2�*�9���i���b^�_s=)�Z����z^ܭ4͢oN���\���zT��*ʹ���
쿈�NRӿ�����\�h�����/
�ꫯ����ﴖ�<;��+��,	�I[��4۹}�y�i72��ɲ">s\20/����~�	�������n�G~�ȍ�t�N���*�¿�G�Y0Z��ot,���K�y�?�X{��׻u����/�ڵ�rNu�l�L�S����X�r�� ���o���_��c�4��;X߸���o��"�3\�cb�	A+,D0bY��,�IٿwW����/���<#a؂��6�%Z$�*�~�И����?
��Y�<�'��7T3ch�ƫ��x��3mB�<X���_u��.R�,e�
�g�x�j��8֥�-1+���3��^�?�x�.�����Ox�bŚFsabE���B��B�%��J���L�dk[sR}�ݾG�K��BŖF+�q�Y){���m���Sݽ�^^����~eE�&`�}�_�ߏS�eyƬk%H*7C�c�Ĺ�/�ܾ��>�ev�y/�����)o��x����������lȊ�ױ�/�>�wı��Ѧ��g>�Y����� �v�����8*���6:Fᬺm߾���o�օ��ZL�����x���������.� ѧ>�)_���]��ψPL��Ŧ������ fHH��8� A�(PX��s��糲U�AHΏb�R���
���:�%���M���D�,T�AX�|��2�D%�
�1)�z��_��_�k/%ſ*PƘ�k-v��Ǫu�kS��
�	$�.a�3D)�9X�Ϫ�C�T�����JaP���_��`!�i��>A�F�!���"��`��H��9�%T�NtL�@5��`�:�t�&.������d��Y�ֱ��ã��̳ٺ�r���2�;STޑ�zŹx�=O����\��x�rX �7q�o��^%��K.��Q�s�)g�`�LN��̵>�����{F��j�k��V��_Gg@�QY����W�CP_p�Ey�⩂~���?�1woQ�E4K9Y0X����Q�෾�-�.��B/�@�@��
D�E��3,y0,BY�
؉��*E	E�D�Q�/����|��F��.=��r�=�C�"����@
�r��'b�,4��7j̑� L@����ΪT�EtI��Z�ipN�s�)���2�J��9�[��*!+[qU�d�c+P��c��cL`�!E�ʶܻ����c���x/�"&҈�(�]p~��'ltx�=���6�kGz�n�[��R�"@#W�<�,�Q돷#�8�cqO'��^zzs�-͗,�93�=�,�'��X����Po��@�-�l1��s�v�w��x��_�m���a�g񙆓���k�X��sN��?�Yͥ��q��/u���d��M�\饎�e�Ъm|j�mݶݾ���x���k4�%0>�Sݙ�����
�J(�E#�x��21�*( b��JP0*-�6�'˓E�LD%)H(]TQ����'�������#��Y"A�� )$��n���V(�eM�_�X�!���w�k�Ϝ��{|���3a�#`e�G�q���C�Q"�N����wz%��x��ށ��4Шp����5�Dzyg�\u}�A�ɱQ+7�WI�F_��+�Y�MU�-�D���X�]J
#c�4�mE��h�s)�/+�s~��l��r�AG�^�L���y��
2�JwH���o�F�G���xR����p���y*s��N�j#���x����e��RT�^�+YU$`d�{˃+�mg�wʭd�!�x��;�g�UC�e�C�^u�U�(O;�4�H���T���&�5r���| )��X�vK�ɢs#���d��'���|*=��Q�?�ѹ7�AX��? �]V��V�zY��k�J�Z�~��`���)� L^������)oa��TyS��UDN�[q<[�?XW*/�h�9��b�sC(���'��@&�kdl���wHA�
*l���E���~4�C�.���%i�٤��[�}W�fΓ���̠R��M���ʜ���{ �v����6��=���J@g>�|�W�*&�{docpѷ� �bzzf�ڱ?y��2�3Y�6=�%�S�!����݋�S{h�sT���g.̸R�t`Z��m�ˈuWD�t�%�_�k�� ���`���`�F<�k`�I������E���'?�Iߔ�A�p��?~-W,�����W�v&�)���,PY���c��|4�N� ת�c���`�^\R�����p�E�YpLE�8�0Q#m�K s�Yo�f��|.�iމw���L#�de%�u��iK��ol�+v�0�N\~=o�yQ�D�7oRק����T�X��x����p�u�0o��$�T�GU,X�s�%�e��X7F��l ��{s[�)7�j�	�d�I�yyh��@溪bB�AmdD�����y}��_�}N�7���������̟�nȐf��J_�&��V�Oϴ�ɣ��~�ûlp(y����ʔ 6��F�$���&K���6Z�"�~�E���f��d��m�z���K�1���R&,����� e! (���O���-n�IH�d��h�h}Ja��#��%oɲT0W�Q�'z�+�:f�"�x�AB���E� �K����0R�N�
��F0�@�R�Q)1
Aל�ZKi)�b&���<������H�a0�7��%�5=	 ֔�y�����l#�1⻕�a�r���I!���g#�-r���X\�ۂ�Ӝ�f�Y�i�%%�%~a�;%t2p}U��t~�Ԫ��!*�8�W^��ɑ<!ŋX׼Ϗg�潒�HX@`��dՍ��'m`{��J�V�Z���I(Zg2L���Қ�� ��}5�x���du��Cm�ܵ,{i��H��Rő4��0�O����[9_p�^��w�>������M�{d�S�c�,�����˳keMŠ��T HG�B��x��rs�Yd[%�D�dh�r܇(�x*׀`'\�d�q�QF��D��7�hΫz4�.bYDG*cy��[FgPS��C}�f�u3�ۿ��΍����s����<+�*q� ����ׯ/�S�]�j��bs
&� �G��<)��R"XΚq6K~OJ��[�E\ks�,b,"Χ��2�ߨ߇ ���N�C�VL��<MQm�3�۩�1���<��|��6F��~��Y�H}���+�$x�PQ��<��QfK���0�־A��\��G^�d��3{�g���y������_,�i*��^|��2�a����^_0L',"�}ڵ�r������z,��c�,LYw�?`���>���x�*� �BP����[��#�&��,J���Hu�`�}�m�y�G�x�l��1"J�P̭�%�n���@���8V����͛zK��,TxO��I�L��Qָ�4t����Cl.�A�~���$�8�g*�=�f#)����ߏP�{E�¸)&#o&��ϕ���܇��R�ϲ���D�p~]��}���o~ӫ���?�q��C?���eĐ��׬C�劯!�F�}��1z����ح�0�j@��EL9��큪�k���/��/�ܲC��h���;d9��Դ���zt�&�F<9v������mL�(j�oh��Q�H���΋�#.f�
��&P�Y׫�$�#g_�X�F�'���{���s&�G���*X-���P�^��+Y[H��!K�&^��Y�xK(�X�ZZ��-?x(O�q*)A^S�G,I0SPV����-Ԑ��<f�S4�͖�"���ͽ���*�`����-'k�Y�y��5���%zp{��kDa��%(��vT�Z�>�`1����6<�*��Zӕ���j�i,k��f2�H���HY��}/�r`F��e){������Y<\�@PDw�!�u^4%ܦg��R�����9GW<ZȲ��Q��b���$���~���K(�]�ML:k��_���;��$�:�[c�}_�sӼ�p��7�SA���@y�E���yw>/A"��WF�^cJTQi���s�j:�֞����4�߹���ӳ�wLcy%�G�n=�z#=���*"��6K�P�-*W�,�w�`�����<:��)���Bs~���x��PL��D�P��zS��s�[ƙ���dzɍ�"�n�1�:iN��|��¿���5���6y�	(հ�ZY<�'�]�/��z����fV�g�D	�J�m1���[�i"�:V,�SP�S��'���}ˊτW5�κ?1o�㗒yH�JTN��,��Y�m����ڟ�=�OV���b���)�d1���O|��1�S<��D�%�y���He��;��G'$ة����^�������b�u�T��'w`b�&Y��$k�{�f]�X_{&y1��z#�1�ǲ� � ��ڂ�<�k��;h>y�R��baC`��@�xn������9�Cc/0�����F/2����,��=���X�¿�m�6��$,�k?:U��m¶թ��6Fw�7c\0b�t
�ο�ń�4�C����F^�������5�f�ĲuQ�IE���_�F+��F�ә{=�,�Ҷ�ע��:b#��<���&�'���a�#�FU�-�!VL�W��(/NTP�(����� ����wu
���9у/L� d��Ne;�!ť� \1��S6����,߱d=[s2��	�	/�W�Z�!�\[�j�-]�̃��t<����.�O��ؒ�����Plѧ�*%�h�id�Ǖ8D��g0t��)���d�������`�9`���E�pl������/{���DV�m鲥>�Ln?cc�6�d���Es���
�B6�Ц-0�N�W>.Ta�L	�t���(�'�vۣIVP�s�⎐N���Y�A�N��Xݓ����+u!GTz��Fe�n��4���M"B�����.��~XX�w8�o�D��9����w���{^ÇzD�b�������\���y]kGA�R��	r�	�ס:R
x�� 
 S���p����jVճ����o��=�P�m�>b�G��i�
��*�G������|Kqʛ�BVv;����$����iLi������u�o$'��%�<1��o��\����y��'-+����ױ�k�n���vZ��	(}�}�km��徙֮]�Ʀ���f��[�~��<-	�G6&�@�տqkK�D���f�p����v�
���`m���i���xq(����"�9"]0ޓ���y�qn�:���v��y�}����O�J�"�M�﨣��F��w�^��~�Cr��,?������sX��\s��7��M��W����_��_�b@���}��zPԮ!�Tɂ�����*�G������5RD��5�C�9+�	��O@�G]޴v��p��,�JF��9y�q���=mKl�r[Z���J��)����$���MO�j=�G=��b?�'Avj�Ɉ,��
�F�q�Y���>���m��?X��%Mf�_�'�hc��?Psh��j7��ױ�?��f7�VGI���s��n^��Wم���d�(�sءk�g��)�'�z�]w�u�%�41��o����o61�෽�mnݱX���/yIg5[S@uY�>_��~�~7!*7�xV��18�4|-v�K���������{ /�	9�����VR�o,�D�����:2	d����C� k-��ɉiMTp�D�Ku�ԴE��=^\$ŦGy�8< 	Ш���5����E����iT��?���(�����n�����.U2�%�Ջ��:5s��U���k�:L�\y�u���-�\��ǾZ��w�@~����,bE|�w��C=���_b�]�^�EJ�ܛo�E��=���v]�����l��n[~��=�ȝ�>�~ g�v��=`䙝Y��$�)u�[�f�x�Ŷ|�R�ԎO��&=�ӯ[Ln��I8�����#�����޸%R����]�S���?���`_��ל��~�Wx!1<	Tc1<R+ƓO>�/�>�����3���ҏ
����	��Q����+�O�����;����R��I ���תe���Tc6���j,��CQ����Vj/����}vֲ���l���:)q<��K(&��}}.*o)J�n���uia=�n��s��݉-��-�J:n~l�^_�)k�WD��9�6�VS���8i����������#��j����'�3��ח��d8��H���E��e�'�,Kط<�E/�K=`�r��V�q71:n�sn�'}�L=�ܳ������m��<kU:yy��zꙶ����C׮�+��F�=��;��IF���>�9��N��3N;���^{��Ǽ\0�T�+����\d*�L��)���,J��~�}��fk6�Q)���
�"I��Ijg�3Z��<�x�#6.n~6�m4Y�p�I�X,�o|cZ���
.��`��Nq�9)g%�}�"svr<���z�Q�����VI����}���I�ޣ3���l\��{t,�4~?�WJ�)�K�)��g�3������͘k�ǈ��ێ��Ȭs�w��y�������q��z������V��hbZ�d�o�fO<�m۲�1�ի��I'��%����)��d���a���g��c�G@{��V���\�d�Vl��ەW��IcjĞM����~b?�$ؓ�54�'|��m����9�BW e,e5ؖŀ�Ǌ�aA�z�E ��&j��I��5im�[^�="_XV�g�Q��6�P;:�Pu2p4�	ୈ�a��4��HG���y�+/A�wI��r(Ы2\ץ��=<)���p_L��1�O�ڪ���;h�e��[bj����b��mt���^�!Gk�!��������M�~��ݓ���^
ts�>^�k^�;��#lb|��Fw�/��~�������l	r&I����y�A;����QGW���w������.��|��>ϑκ�c�+u����Sq���g����u62�ê��my��$䟱�]f}G��� ��:"�w�����9�W��J������g�E��br�>��F����{�x���}���*���;�Y����k�+�$'a��6T�+6c���덂Q���*9��-��_��L�+����P�G���"��9aD�"���1^2�2���|�
�1��n���(���X]���2�w�����GM}�za�0x�r���w��&���3s���gG)q�?�"Y�q._����*▍���g�d)_�k�8��f N�y�+_�kO_y����?�coV�o�Ϳ�?��?񹈙����?:6l����Ϟ��H��#���Y�i�9�A�뮿�N=�,;�����Î�N8�6w��	!���;ow�!����j'�t����X5�?��F[�jȎ?�����4�c��J�W�1۾c��%�Ɗ�k�a"�ُ% ������C�1���C#0\�ˢo�34]��t�c�AZm']��Ϊ����<*���������Z�^fA�H����6��"]K�������X�y	��>/ap����e0ڨ�
}�=�s�;���E��k@��;�����;�)ԧ e��4's����#C�f�3	o�S�����\�����^c��#���:�,�����!u�t�MN � 6��u~�9�V�f?l�=ro�)[�n��?��F�G}O��Q����ϭ6<2a?���X�'�֭q"
��=�Yi�y�^��X��d��v�y��iR[^5���n�7��r[��{k���"ob�N�ɢ�8E�Jε���<xKa-�9����*ңW�EQ,7���p8a�ެ��Xp���ٽ�����}s�M0:��3����R@ΌH���Y݆�U��N�������)�/�P���ΊMlP�*��y��*�8��ň���ǡ��ӈ5�E��#�TВ�'�C��b{	�={�uf
 �N9[ڿ�S$�u�?�;�:����)��X�|'xM`�[�pσܗd�2[�z�M���FQ�u/�����a�Q�u�s���`��w�{lx���v���E�����w!\��g�ޘ��ݝ}�����NZ���`j4�=Ѣ\��-O=h#o��/��{׻��X�� Y X}�����z�j�k�GKMp��ǋ�'��%�c�_���V6�h�6#ŲS�+�+�!�XL���*�|����U�}a����0��RL���k�+Ll�Q�C
4�q%�s!.
���	�+r�9��I	h�u����B�뭲[�e{aÜ�q��}W_}�{��f���|�����ݣړ!�9�{��s�l������MM&�0>�{a��¬zg9���z��f��
�x¿xT{�����{��ղK�V��*�_�����¤���P�ȳ--���
�����eu���{�m_�e��K� "mADE�b�h���-&Q�����"��b�-�`��BD�FT�" ҋtv�������|��~�9��{������ܳ\�ַ>�yN���]�AY�x��%/	��������,���k��qՒQ�>N-��U.���f��Y�x-C�(N��9>�#_%��lk���bm�m��R�f}e=�l��g]D�)t��8�����|�]���g��X���/�:�|�Qh))JUH���<ήJz�ĸ�X��u v�׫�<某��c`YW��؅�[#��i�9~:xp�VdG�.}� �>�>ѧh>*l�e�;4`sk��q8�}����Ͻ�֮���2d���� ���zu)^���oV�':0X�n�`X�|��$�H1�É- �r����� �F-6��A�bn�\~�_X��$6�`}��Q֐�?Gǘ�^i�öYub[�2�═��Aơ8h 9.�Hʿ��|�X� (�FP�V��H|��{�j"��~А~���x���V����7|ܾ�8tͲB.tL�`g<LQ5�L��;5�,���h#[�<�s��ʿ���a��Yk�=eH���\�(��?�nr�c�Q�hw��.ŕyvg�5�7l�Du�n$���Y�/�"�����X��<�Jޑ�nl���۲�J�2�eO��)���wo���w�)ny6]�W�8�)���1�0��+R�ʩ�|�{ʽ)�#���I��O���]�7{�����E�Ѣ^5R7�L2X��e�s��$�|�IV���Qԋ�o�L{�4��e�����ްt�n�)8���kV?֬Ò�W�9�^����%�Cm�3<��6������������@ ^�e�h�Ǡ���/FȂV�2mi�T�b�J���bT�H@_!�H�Gh��RӾ&J|XM�Q�y�b�",�u���.�-PW�����`R����V=�Hx�I���Q9/���JX�t����[n�3t��y�Q�T��r�%��:�[�떱��X�^�[���7|���8&�tW�.�v�����~�oX*ЬZ��/n����Ï�vTN����7��Ƴ8w�q9}��3Xy�ќ�MqKK�e	ζ�egY��|$P���լ<��I��S��OsǗ�����>'*��������|�0��.�̌=��>��]tQd�6�o��݌qu���¦�=Hݑ��m Ϙ����;<�ȣ����]����"�2�z�O�4 |7��J�և��7G��~�3�mrg��w���M�{�N��`�5{n8ꨧ���=.,^�gN?@?OY���s����Y��E�j����7�y��=�4)ShK[���p����(#�Q�=��l�Դ--,�5����WD�8�a����m�<(�����%��P;$��u�3CT/a�=��fox������j�8��#�	+��:�ظ�u����?����R��"��dfZ��&an
��/*�+���85�}��ap�?�ߡa���	kW�
�7�7��yX򥳣'�^Eϓ*K�����0��2@��Q�*���}p{P�L�|M��a��2��4�k�TO��C�7����a�\���e3�o�6jz��Z���`�	ƭ�>V?�"���+W�Pm>�⇹_���I"�s�!����懧���s@��Ca�ڧ,��v�,�=�[�(���Y�B�7�䧡�ws�M�Im�����vا(��	�	��VC�˾���j�S��SN��˼��¬��aϐ��VK�x��|�;V��V���e��x��h�nv�@�ɏ~�c��a��Z�CP(�n��۲������M-��q}�-ʈ�K�N{�*�s�����{J��n��p�Yg����}�d��#�/E_@��
B'�+�/�z
�^t�������9+,�u�%�}�'�,�������_�첼��r$�-���E^�&���/̒QI5m���L����ζm蝑Z-�6eE_�r�e�a�k�+,_��W��>��O�M��T+�_��B��@��mT+����g>q�rN����ծ[���%�r���4�<��wɋhDR+	kO�,KO	6_il�`����%?��U�V@�?0ʒ�_.�x�ڟ���U��:0����y�v���(9��Q��Ch����E����?/��� ~��*DЧ0�{(���;�x���g��Hݠ}P��_�����|.�J�'�]ͳnf �:�R9>~�!�ED�o�`�P��}����eM��R��c}�N��4���~�㟲���^�|O��Ю���#��!%)k��MB��e,K��O�h\�"b��7�#̂��0�ꈕ�+6=d+
�}��TV�k�b-�����yN�f��G��U����
A���3���n+�&������O����?G_d�Ϫ�):��/���i2E�U��v�IR����i���f� �{O-"cf"�r�?�A]�=B�_��W�k����eFY�E�<?��,3\{�V�s��#?��T����f,�_�Ѷ����0��=���n��PTG���R��&��o��P7�6����yG��޻�W��+��s��i�Q��C�AT�°H	8 7S��$�E� ��J���ۙ%�dmx�6��-B@=�M~OG��X4"
�RĈ&����j�,OO�e�����h'���.ޞ"[���5LjI�GA����������&MGƃ����i���2N��E�k3kV�Q�Jɐ+i�r�r����W��($�y��mA96%w5�՜E0l��/�B�&�\��%�7���1�ph��~sK�H�:���>k�H>Č��j3�ᶞ��?U��9�����P����z:�j)q[�,�tp*$ �k�z�ue�{��&Fb�t��(�d7���<�y ��+�q�WGY�ry}�F��� =7�?��s��t��X��u�v�U#j
�� F�LDj���m�r����H,
o(t�SnO���UDcK�Y�'B҈:z2E���;�1����KII���@eT�o�q$�~�9�OCh5Q�0�<�@��H��QJ�s�/H�[� ���/�c�h/U�(s����z���������>���)���
���>M8;\Q�&WR�,��lT϶�,�� �b���k!�|�;��c-fċ��ѷ����',E��1���[�Z�|!J���X�s.B�t=4h�Y�:&Ÿ5���h��=T�������Gu�X�;���Sr���)���=S�xD�!�U�Y�IcE`_M>٢1�á$;���б+��ΈC��ԒQ�D��'��W�u�Um��)<�n~1��8 y�˅�Ȱ5��f�%BX%#�K�~���=X�J
�n��M��Dj��V�K�����?KWm�MT6��ь��U]����\��)�	�w�+m͗)�Q4ΙE^�p˾� �$at�W�}*iE�h{���qkI=e"��m&
/�2%�\��EMqT�Y+�;�[�PQ�Mݴ��L�z(sQR+�9ޘ��-诮k�/�m1f+�w���dS6{oᘸ�,TB� >�篙Oו,�&o��y�	�Q(��s��)�Сs�O�_����2gNOn�#D4��Bm7k#y4XN�Q�/��C�1�a�V�6h��e_�J=�7��Zr1�0)%P+��>?���)�jV�7W7��7V�Z�u����4T���|����{�M��=��1��n6�=)"OC�WT�Ÿ���0��l-�E*/�,�re�v�0٬ �os��$����>,�d<��Aw����U�E/�!�@��C��X ���/}I�m��ro��]}��Vs���dJ=��Ʈ���/�xw�dd�"R� �'bl���$2BX��x��DSH/��-�7.�o{z�,�P�s�m�W�(�]�R��!:�d�y%M�p�J�J0d��\�aK�A�����~�s��y=���<�տ�Y����@۰c��3���Ot	B<Ǹ$�c��p��Q����b�����n��-��1�T4��șlM�k�B8�evi�x|�+��T��RMR�w���B�#d��q�$�uHť�b}�"�h���Ȫ'�@� cJ�ʾA���d��>~��*̼�9����5�8���d+���IG�*�5�&���Ƣ΅��k1�$�ܟGQ|��������x�5؂8,�Kc0����馪[ �a�m
LʉU�1G;;���\(��P�\�|LZ���u�!�ƿ���Q)���l
AC��\JW쁡T)��;�)r�W.���(&��A��H�=�C���{p4����h������g<>��̍�&��8Z� P��j��eU�I�s
x9��;��H���9)t)r>�&�硲*���#
=�O���X�"ߏ���T�E&[��ĸ�CD��*��h�Z��
z��-T�̪/%#�Gڽ� 3J5����ǩ=V	��~��&��[����\�W�Q�y������5)Z��������aJ�T����E8��Uμkiv���~���7�@�����J��9�ƴ;�o+2��x�::+Yf�ìl� pߌ�;k� 7Tqq���F��7B?�Z#񿑞�ږb�����|%<^��5�h �M*���B�c�R��������H��EM��\�{�"�7����;�;O���;�֌R:;���x�o��!����iҎ����g�C���Pv�Vݛ��g���c��E�wnM�y0�chA�}�g&�����3W�N���ם����`�ީea+Bf�yXI5A}}t��2�s<a�i�����z�IM�3���L)[��m�H�T�)e0�5��"@
E�SL�m�_�BXF%�)�k�c��L��SD~x��d'���O�z�a���m"��V�7c�X�_罴����}K��z'��|��exoK�TA��[�mlb�ް��'=J�x�޷���ֽ�tY�=5��\�3�֊�(?'u���|�ӣ������ȡ�S��Q��T�F������Z�q�CU�$��y�Y3iy�!����o��Ψ����)nx޼���a�:KΤ��(aҹ����M��h�7JVB,������ ��/Z�>f_T�� ��%哽�8�9mmry[$O��J9W�G��U�x��=�x��<9-�x
1�Z��S�L�xX�{=�Z��S��)q�v��&)�V�I����"Aj�a���[�$)%�v��a���c�h1U�I�� 2\��&��h�VO�q�Q����PV璵��r��y����s-,M(��`s�V����:`�A�����,�ߕ�����p�QG��sS8]�\J�}~}˯��<��Us"J@M�y��3��{��lq Aʊ��_n0Pߔ��58<���@�b_֢�W96S`�|����~���� te�q}szYt�WŅu��3���
!�d���������d���־��V�1�R��� �c?��f�7���crkI��b���?����j�	��� �[��ih�/������B�Y/*����ہh��K)�)��;��}�1F�ĢE�æMBGg�l�y����52+J�X�K��a��/^b<�rw�m�d�v�a�����y�T�9�~��������o;��W�J��q���w���ۢ�"��|ޚ�R����)Z��f��Dy���yL�"�u�$W�����.Y��&�S<~"��H�z�/U���@D?,�e����{P��M��D����8/�4�y`��+�YN�o-��A��-��Uua7�l���x}QS�1T�e���3�����~�Zu+�
�y���c�1Ѐ�)��y�q����~��[r��$U/'�iXq�I3��Be�%K��A� ���AR��eɀ%{W�^c݆@[tvw�=�\�X�$�_0�������������{��^'�/pMn��_�j���Q"�R���/���(���b���=yWq���B�ޢ-�#��믿>�
����B0���U���+o#���xg��Gl�	��ҡb\�;�L��E��Uա��>g�y�s��1�W���>�_g�>���=��¶���q��?�����=蛡t J�����'>�<Q�y�E(���;#r���[��H�QI�D�澰ے]ü�¢Ż�����ʹw���R��k��^������J�ț^��4gx�s�-�y�TNK�~�âӢ��O{z�k�ea���V���f��C�A��.}<�ce��DV���6@��XZE_T~>\����mg�Z����?�c�¾Ta-*
�;-@=	r�P���*>?��#I4&fb��6�B�\���?F=lUU�f[%��,a τ���%����w-(|?��s�T�2?-����u��`h�m?~_%�Ѝ�������*��g?ks�¿׾���P�P?|򓟴�#T�ƴy<���#?�@'��=em��֭��"�i���Jٶɼ��l�΄�ǳ�O{��L�ɝ�g\�l�p�����&�|�/¯o��ݐY�������=�����p��Ǆ�p��X �|�t�bWEA�k���lٲ|" �JV�౎���'��mU�H�6����,l!���F��b�ɡ��呕�a��}�"=��������~-�o��|��0ط9��prȰ��Hj!-yL!��rHߏvr�c���g�����և/~����LY11��ΒmC���ů;���SO��:8���^���/��b[���7m;�9A�������@�>��G�7�����'���=��~����"�(�:!�C����|{z�V�a3^�w���`�شV���n��e(*�êU����-���a��e��]�f]�ߟ�8�\�.�}�����'[G/�w`аYYY����c� c(yؖ�+R��OwԶ�jR�*#�oB��;�p��z*�4�)������p%+�V�U#�z)q��0̖����]��C��ې0�1E8������'yY\~�������ֳ#�0.ޠ8���z�E
LCu0��ۻ�=��*�a�����Ɯ���S�ׇ˿�p�	��7d�'�n���p�]wY$b[��i���&E^p�E݃��|�����/¼��a߽w���#a��}��b��֮[���p�?	���ߔ; �fbrr� u#�+ĀO�]A�����}�(i+�)-�e���"�C�������~7S�s�N�<GOs`CV��5� �~��hd%��Y��?I�Y�U[J�Bt�kr/��HG;�C�����cm���߹"�wιa����&Z�ᔓ�̛֬~*=�x�4*UxҊ������Q�$�a��Y��:�?@+�p��>�W?�fU�я�.�=��2�p���L{�J�#~��K��i�{`s_�;�ۚ*<�όx~ظ�'fq�rW6[l���u�6G��Gm�?�\A|��Y�SLX�
��'b5!�|�H[��-�l��hY�SY��y� ��X�a�0�ը���8��Ba%��b)U�fϙ�'�ߓ~/.���^EV�x�V@�/�
�^w�u����N���뫮���,���^>���Q � @��#�S.U��o�i�c�°�^KB��ު1 ���\w��`X�p~����-w�{����@B�ΪUOm�M{�_
�M��;��sٞH�C�#��0��qY�������\�a[X�<'	,�/��~�����;��=��!1��f1`��җ�d��3�I�D�ôe��p�J��h��^1׎DB5�bHJJ9�laӭtf�
��BZJ-yC1Z�n� �؜ΰ��Ѝ�T��I� ã�?���B<��Wq!�hFZ���O��-���7�l�n�Wy�w2�V�ZV=�xX�����t��l������T�2n�Zm�E@����L/�0����c�3Ꙕ��p�7K����ņu�CgY��MiqqʤV�6��$q�2B����� |F#x��|�.����t5e����
�Lm�W}�#CuYM�=�C<��"�r�`dl4./�åa�XH͈ޔ�5\F\ �� �M
?QØ�@�P�ƅa|��;�y^�2��z����s�����/��'�c��) Taz�CwO�u�d΍%�nI�4�
�Sփv�k�L���o&)?�4������Z���S���:-�M���v�OWGw�<0��ss�ӀQӖ����4/ݼ�+�s�9���~`�_����芧��֖����K�no�<�4�b����Q��r<�h�1��D�G?6[�5*�ٶ��u;O2�>)e��Z�	`��::��M�_砤����@;���Ë��E���/�x��q$��k���4�+c �Q��e �}�O<�.�E�ڊ�Aӿ�=��Pn�R����`G+{����ʺ6̟7� Vs,�?��tǬ8@;�������M�;��I� �"�Í�"O��$�2 (���#�?���?��?�/|����W��/(���-����S��{�.���6<)Z�C����V��k�eo��������'�������2ۢ�j��;j/(+%��E��*tQ�y���z.�����WCw>#�G���X?ߡ0�a�
ݺ��tu϶�J�fx�����5{j����ua�^;�6�gI���%�R���C女p���+��nV)u�q�psX�vSXs�TI����6�n��=b7�?�b�<n��ִR����t���Ȩ�;�n�.��_�o�}�C��N+\$���e�cnˎ�ɄZ'�TQ���(i��0	�t'�P����ڐ%q��*Y��?�i��xF���O	��`t!�d@���.� Ý$Y�_=Ҝ��-�fT�:�֦�����a}X�~]� \�g����x��C��Y��N4 ���MF�F����	�6�
�V�����{-�#���;�7���W�5�����Īա��k���ƀ�����B[�]K�i��s��VD���p�aO��zsX�a��*����[騄����~����ͻ��s�N$ox�����jx �@l����g�"�EEBB���Ԗ����5/یs�_u���������uM��RW��U�P5mi���j�����\��_���Z�v���-�V�%�<1�j�ق�!v�����I�U��9�<]�O�����{�Wx�oSX�iM6�g���U�[I�ݬ�粽�I���Z>�߰1�u�=F):���d�S�eȚ>몃�?�C³�����Ǎ��'J����3kd8����Z��QO;&�Ǟ����k�F����mA�g=�n����j� H�PZ~���t����-h�Xpmi˶�o���� ��w������y}���z���ʯ���Q;{�_�|��&(o�=*��>�ݴ�8��_g��W(��ܠR��\H��/|���^�2��R�c]�$1��0�|�~��������t���/<����xU2~��v[N{�s��
s�.�c�����]w�6�t��;c��5���T��!�w�WZL~Y\�I�{���|�>�Ʀ��G2g��ea>���ub ��e�p�~���VOa��
�ָ}(�W���:5ߞ�(�����J_O�M7�d�1ա����(��� ���O�H� Ҿ���U��J�����i��R�导� ��9�=�г�q�f�!`���A�0���9>u���W_}u�m�Ea�ys��y���f͞V�z2��m�r���|�5����7��^{ì�9���U���o&iB'����������a�����a��9T�����oF��~�j��FTra@��+v��;��U�<h-�do[vv���
w�[U���o����r����zܨ��0~r�?U��ߛ]�z3�f����z�*�J[7��,���
�b���׿��]�O����(~y@ZL��^~��-�=k^\ ������@�ي�2cq���QGt�u��{��U+-<T�3��m���q���Zޘ�%��/~�?����7�����q��W��6���ׄ��+�巈���������fx���;�>������28���w;�Iy[ڲ�ģ{<���jCi�ݼӮ����m�$���y��6��gaTY\
`Ͱ��l;�W!��"�c~����I'�d�Y��	�b�Q�N��������O<eq'|�;��:t�;(b�i����On��y����S��*�^�7+�R���m��fϝg�W^n�����u���LY6i��?��n�:(-'��!]$�����>����f�q �/\`!{�ψ~�c3,0a _�5=`۲}e���L(��̘������@�u�E��8\�`��vBj�S�UΊW;�ݲc2�Y��r�c�D2t-~��`��>I���_���l���MA'9�o|�F��^Q徘z�B����|�*�n8萃��˖[�?�G'<��#�E`4��\�6ܗ�3�B 0s;y5asey�jg�ǒ������X7��?�x6,2���B�=����W�j�\F�O����
�����G\�mi��*��0��ϕ���	[�V����%�����{.F���O�f��Y�[��A�VT��OA�5x.�³4jBA���O�~�к�{�F� �
���Y���Z����O�G{4k��:+{h�����z���xB�X��}��]�5�`-tf�a�q�ש�Q�d
��J�!i�!�Ց���^X��/�� $9������e��V��(`[L�V�}�X�FZ��w~K�@�������	g!�<��/�	���5�暩�����:�*�B*���{�"X`% ���~};P��HH�}�mn{J����3�Z�V���Xv���ζR��Ŏ�ي%tS��
QV�(�T�b�'�ݡLq��ϊ���H�ߏ�C�{�Ï~�#�ü'����J~r�$����c�CF]�і��7��V�e��vU�F_�P��J�⌝�ʟ�݄m�TMNu�g�k�E�Ɓj^,}�9��L>�z�<H� ���FZ����7�).&c	�X�WyAS]�#XQ"Ucb�
y�y����C��Ct���#�+.�;)�c�>����[�o�_�}*Y�R�o���']F���X�ԓRP� ��^��͏J�¼s�k&�jod �����_�����Ð�}��`��<PO~+䞌�����1�כ�(���?.���Qyc��^ײ�6�^:9�܅b�@�(�z�[�j. �[�����e kLx`�f���N-uo(k/5nbK-�$�G�=��A�K��N�Q��{:�f�Ų�EQߓ�>
j½p�[XB��Z�@-�gX���u����MI���/�B��g����D�@��(} �]�V��9
�3���[���;��1���p4t�J6�E��E#��5��(es"d��>q�_#��j_�̜a�R���w�{T�W�͇?�a3�t}8jd���Y]-;���%���]u��M���p��W�(� ��|��A�í�x}(��hpȂm������0�({�Ϛ*�r�?�V�T/2S�FEp(D�b��𚸈��=^�Π��E��<(zAh�e�6F)�d|�����I����ڱ�A�����D�_�GJʟ��$eP��@%>(�8I��WD��͵���ͱO��fVO��V�Ŗ�R�fd�o�3�<7]SY����~�%�Y#�Zy`<��m��fc�^��k�u� MhgFf��yK��rke�+�Z��/^�r�/p��`<��ۥp�&D�%$&?�#�`��R@^���5�e�*l#��lb���>�*�U�Vc��-�֥ב��B�d��R<\JQ������^�F~�����Pl&/y##0�P��țsF�)l%Ũb*?~�@d���K�Y�v���&��l��ª����Q�@�t�t�b��+Ua������Gख़��gˀVV��f4��6���暊��z���sm��3����tq��W����V�~������R����uq6?��=��?�IG�&-����($��m6)E'%���>�z�>�.Z1�k��&G&�X�:�֑Gi
��@��>���}�/�]�\�ue1s��7�Z>���H����
e"�N�FU���0$����jH�Q��������1L��������<\�7m���I+��c�!/Y��pH�o���?��&a;o4H�3��a~�9�;ƒ�����FyzJ��#-*�Qa��s�O2q�~��W�IǺ�z/r~c�(H�,�}�))�)��G!yإ�<gx+�_�c�X0��؄��,�~eD��M�䔬���I�s\�dI�O�gAn��Ip>'�A�)�t=��gk������,�f��ZȔpTX��%�s���t�:�9'�!#�EC��z�#�����M�K?#�~�;JF�2589�]���,5lJY���Y�w���04�.�T��0����tTlQiz�uBz���jg�j���9���t�VR�Q��ku��ʴW���8�}�Qc}�V�����z)g%"�KO�UB���C�DV"x��+7����?
DI-����1��krj�q�b3-R��z�rC��5cA=K�ԑ͔��x:&ŏ9V�[H$��PD
1�D6��;j(�筧�{�~GAWh��=��A#��b]K���Q��(�;�<�&���`S�V�J�S�HcEH1�-���܄�Ac��W3=�~kԱ��fe�Q{���к�J3�߬·R�j8�a��ڪZ�IȔ��:-'O-B�db�zG�k�'��/�������ڷ��5����J $q$pa3��w��h��0)�=��::Owg���j�����5l�^i������2���#-*����^�h�q_�&���r�0���=e�g�CǪ�i���PЊ�9��E��YH�63^�o�;
����N��!;ϸpu���?d�,�t)�Q����@H�{�+]'��3؊95��0VA&Ǖ�sOZxձ/�0�E�;�.�nʍCc
�:�s�OǤ�u4�Oc��i���a�&�c��]w5*VU�z��Q�d78M�=Q�����h&��w���o�a��e��
ӣo�(�&�b�<� դUa����)�YY8R�,��$��ީ�gx,�����'/O�s&�
�
!�R&��QQ�����ߔ���(�z����^�+��<�Ƃ��p��<U�1�h|)�%e��������RE�'#�X��?�C���?olճ�uZ���e�]L���	՟�Z�9�:�����PP�'�Y{�4��	a�Y�������?�䨄>Jm�:ʝ��m7?���OJ��P�E���_V�x�]`�KC(�j۷y �}Κ+� �u)b �� �_~y>0&�:�.�&.�L���g6Pe�kA�v���,]���j�l����W������=TL�
�M�ܟJ�'�T�7�wW3"��b�0c�q�x� Y�Eԙ�c�#)�E~"D	LY���9yT�Dqr���sնx�׻���TG)�V��/��\�Ej�:�K.&x՛�!5M<G
�)�$���+�cW��y�ᤓV�=��==�J�7�m��Px�Ǭ����z�Ø�[XX�ɴW����]mC��3�8I����n����M�q5N3�==i,��U�BϬ��Y0���B~<�I�l 3�T ��&���Am1L\���Kp�f	[m_1��!��������O����b�^� �$��$/�Rca*����(�K�$����Q���E�(�F���R�0�S߂r�a(D! ~ON��2d���z�������﫝sJ�Y��XT���t����W�e1���{x�P��T���q���q$I��!r%[�jIX�d���z�<��p��ׇ+���NW7׫�<i���6��M���I$��N%��o�J]�d
��|����c��@�%�l�ޡo0~?��B�pË��v����D�&�?� Y%*�A��'� ��K���	ca���<|t��欣����u��ӻ�
oy�xkE@�[T� �(j��7����t|��b"EJU�A��X���D�U9	��(��Έ3�3�󂹧0k��TU,�w�qǍ���ʯ+4+��T��74&tnԃ��cn��؇�FOPV�+����ܳ�	'�8!�KI�˥Z��;�d|��q� �6�<�0�<��ʧV�cc[e(�ZCӗ��l	��>��/�ma��w�yG���_��}40�
;����V���?�~'R'7����&�,f�;�!�� 4lrtt�A�i�X"�e�w�.U�
��f�2�����lU�����
1�z
��(>�������M��SY�:&�z�F��>Wa+�����1I�,��_���S&�x!�B�SS�õ������4��&�����3��R��������[��ݏ?.|>��`���o��d�bU��v�iv�4����(s�'�|bڏ ����3���w�֬[�ſ|��ê'�O{�3�ҥ�����-^�]���Ӱnh��e�Z�%cc[�|�֝^�����љ��
+W=���DK�?t�l�bQG�7�p����Uk�QO?6��*�R����N-�<
Y�~Mz�bXF`�{sT���#耱EO�J�AU����G;,|�<����ĳ��8��"R��{x��d�VP�����E���d��ZBQk��W��ZBaފU�x�V�.��'�=m��&�E�|\��Y�F��ys�KKR/�m�������4W��|������}O���Ҽ	����V\��`Q�oi�R����/�{��a]T��w���9,�M}����~���p֙���S�@����([�ʴW��	@1���Ι3;U{�o��M��H�Kw�����?�)~��.�����}���?��!y��7c���z�^hȋO�y6YXF>��cͶ���#4�X4X��,⛅��
p�F�E*O�;ؤ�*\�7��d�Bl���a��yy��M+�UQ�D���J�
�H����"b!-g̞�{�y�Ɵ �����֬��p�C�5��r�~<�Z>^}������o��C�f_��O��p��[N�s�?�lI����
룞Y����_�bx�E�	wYl��#;2<�Уa<-�g���	tW��K���m
s�v�[n�U8���򽉟�5k��;	����as���zVX�nc�����z4�<� m!�x�	<4yx�^`�#{�'�MdYy���������O����C 5Ƚ2���h�d����^���tN�!:��]�"_Q1Vު�ڑ�$�����mC�WJ�U�L3�7�"2�\|ިH���0��[woC�	��d[9~�ܥ�{�dk���И���?�"�EO��^t���1�c98�F�0�U�m֪᷿�9��	a���>4d���ӈ���V�z<>�V>��z�r곭Q�A~�ӛ��F��Z�.ȴW�I#��RͲ�W���3<�أ)�H�ue-�Y��G��ąN�E �o����`g�y���TSx�'���/�5�җ�4��_�e���'ێ�j)�V�r�-,N��aq��M=�d[�SY|�{�e��D��?��Qdx����˛$L���ӱN� y���i�B����~���r�O<�8��
�%��@�+W��{�p��ˣ�9/.��3�� J�[�TaRl�J��<��,���.��#�?��p+���W���PO�B�ء,�����!+��������>��+Z!�ërχ|'�/I,P
,x~G�׿��f	(^���b���M�����+c���V8g\e�QԬF��9��'ק��L�թ��D�PR
��o�C���y
)��~����/.J��0�"O�WI+<Hn���%��+����}���Q�j�ĸ�GT��
�R�3�W:�EtpB�8�fu�����A�E���<�#�^����jQV�j�u��7����՟X�]�ܙ%]C�����qM�:�8�,wA=>a���ĘZ���7B�8U*�jB�4�!w+�˒Ŝ#�gC6�ERS=��E
��'baf,���~�|�m��62
�Qb#�0��&Y���IǦ� ���檼`<\B?��Q���+�'�=x-�a����\\l���e���`^w�Q���OL�uk���W��ು�ƥ����[ݳ���`�YJ%�!�^*u�M*UR^n"�{!atS�^���O��2�L�>�{���y��U�F�8�BGE�f�E���L�\�ĥ3�K^���O~Ұ� '�˼=e�A߶�GDʟP�^O���Cё����~fFA��B񵒱�C@�`
���G�&��	'�`s[ʜE�ӷ�������T�������ƅ�V6�r�_�V`��j�~{��.:�3�#
�&���L�z&}�tRp�kf�ww͊�¡��Fk}m�Y��h�f�QBgX�;�Ǯ�W���?�'}�Ї>d�>&(�?x j�۫ց�(�y*%�&+b4T!�K�[U�;j�E�����F��-*��)  �G90U$���J�W�J�z��b�Ó��]:v��!� ����Kx�0F�(:'e����9�ȧ���k��5���:u�9���u����-�bŊlA������UO�L3���	�j��O��]ʉ�3���{Pxr�C��G�aH��*�P����[������ ���Zgq�f�q��)��(8٧>��N)@�>	5��2��l'%(�O�xK��
�R[;�0QhB2�^�>�-��4��c,����\�\�o��2�h�񊮗�E4J���Q�V�}��P��u��4�p��>���'<��á .��]�E	�gO���ݢ�K�,��E��v0b^H��<M9"�T�_ٴW����#��}�s^�={��5�+,�.�~���~���Ҙyq�8���1ǝ:����V�V���
_��YU	"ڽa񫠊���<jH��2A�Of�_��2�t�bX�8����w�(�;��d�c�|��4变r���ɂ��fAP������@�I�&���������������}����k3 i;��cC�^{Z���ݖ��_���0ؿٸ�6m���ts�qǞ�v�3��p��	�@J��3*�g.�O�2��:+�B��������0{ޢ��!G�E��m�;V\n�.w5���h�@�I%7���d ��ӟ��n�����  ~� Ą(E�KJ����SF䕨���b�0����D������־�4�CV�����lq��
������A�|�q��L���D�w���	>=���¼{e��KϷ@�v���s��>Av��n
#z�~���1��%���·{ "��>!���Q�0>��������]w�i�Ϳ��?��N�,�T�` 1�1��$�İ/`�%M���G��M�
!�k�C�3�f|݊���wb��Sqt�d��zvO�O�����X��w��k�i�j�A%��aNT��.�?�x��E�=w���:��|�!)d��6n�W�ϕ�_c��]��{+3��O����K�f4��=[��Z3����h�����E�ȨU5��j�0�:���M�!\pAx��^��o�&\q��k_��YLLmW1Q�&k�S�>b�����K�"��k&n9^xb�hdbiۂ��կ!��j���I�ce��NQ��s£)�*�@�d#��+�b��c���$�}G�yOD��"+��'���WwM�P�B��E�+��B�B/�h��_�<�����@B8��������E�r�,
R�x�į/�����;�1�c����)��H�D�9�1����s���crO�f��o��`*����d�׊sa?P��M����4��/_ȋQ�󊗽܎o�Ż�9s���?$<s�)mC��>�9�P� І�%���)4�zjB)#�O�z֩,J�:_է�7��$(�!_@�]Y)bGT�NJ�6��`�Il����@r���>` ��\��p�r����0Y�-�˕U�;߃�.J��	Cų��H������{r�RZ:�S�B�Hd=QX��/R�οނQ�.�G�����ENVe=���}�zh��q0V�@*���+�}��Z�@,[�0�}�7�*c���£�������LfOx�P|��zECq�T�KIm�k�����~��_<�@;g#|G�~�Be��wA{H���CW�f�q.ox��E�C,<���/�\�1(P� ��K�~��~z8ꨣ�;Jx~)^3���/䞆�Ȍ%v�����WX��z�M7�
#i<ł��Z!��TYV�D����o?+�Fi��]v�e�\�w���h'E�+\�5�Ӕ2�I�q�9�+_��m˔t�:�!0�Aqބ��;����;L���t0�\�Rǣ�g�{˓�c����(���̹�]����X���z0Cmϓ�),e�C2��T u���gE��!U\ �u(�(�;�qSj-����3�Q��\s���/Xؾ�	�
�"�f������?�+Xy8@�Qp֭���	�O���Y �sl?ߕ{�x�o����g���O�$�'bM�}��,,X�Z��6�	p��싱��x���x򋱮�t��w,:��X���g�5C�Z��`�q=�y��F��Ɍ�zZ�Dq�
kEn�o�"�M��h���{��)��b|>
�N�@�L�`Q��m-��@�M���w�-&���x�O~�܂`���/�{�7V>��$

YҜ��d�� N��eeyŞW �}Ja).�܃����X����+9=�2Tx̋�ڢR��)T��o��d�_�t>~�-��Ň�t>�影Qצ�IP¬�Q��΢ �C]W�	{0�x-CB�E�Oޯ���<y}�7�a#o��Ʊ�m��x��[����2�ѥ������m�$�6ʱ��x ��?����{��^{�:�	�1�(��A�����9�ЖI����3~�G��c�'���C�EI=]\YA
mx������c4W	J���X�X*��b�a��O֤� S[;3�G�_)|3�'��%��%7ٷ{�y��XM����x��5X��GǨ��rqY[���4pM��G�z���U�P�6R�XO�c��ݓ+(�O��ׄ�qY�+�~�H<��,:)1�g���|2��̞~z,eQ�#��Z�-�~z����w��[�K
VcH��C�}���3�SCH��@ʠ�exCL9,>c�1t�����Ka�H}��G�t���9/�/0w��_��WٱC�v����X5�}N�/�X�bDe[\C�O��P�)%��6�><���ذO�q���|#����nAt�"�|q�@#%��.��P��J�MF�Y�?ɋ�d�MB���)��OhY%rk-ќQ:�[ ��z�%�BԾ��P-Z]�da!����?�SM���J����$X9f�l�� ���D0� ��x+�uU��{����Qܗ����a����l�+FΟI�dS�h��'Q�,��(/ΗEoO�J�EPJSR/���ל}���kxl��d趾��ay�׍k�}��5��uQ�����cD6�[J����!$��'�M
�Ѥh�țf�a5��߶��·	������K1yY�7�ٟ���;�7\3§�w>������w�Q��uև�Y�Q�Ωt�s�y7{�\�� �cp6�z��a�&��\`o�!B�ԋ��X�B<�#�G��� D���`>~�d�,���QP�E
PP7<�I>a+/AJD������}�Rg�qFn��!��J�Q���cb`��!�K����-������^JL��(Y�LL��e>���d��Zם�1�u�@��mOׁk&��~�m���|�3��/6����d
�Ca��C�0Iz^{@?�|���X
�#�|e�)<H�k�H8��
s� ���J����'��SO=�ƙ��
E�K��s���k���4�4�=�*���xd�(SZ�8O�����d�)��v�NT��%ijOpj��a�>8G��]�앰ւ�ךk���n@縵R��8�������U6�����2R�>��x���b� �()[M\�A9�*B2%KE�X�P���ؒU?9�ө���R*��� U3���ۿ5�Id�*�^�W���T��hC	̕���Q����(��4[�t<��|�+��ҹj��9�""h2E��#�J�^0J��9�z�ߏMY��������gD^'���'>a'��v�(k�G��vAa�X\r�%f�{�[�iy��7���"��BCR��X�}D<�Ya%b�,:��\�����{!EM��d29��H$�-��_�a'?������Y����Lsр&~��镧���y<dybrJ��5p������Ʊ�� ���#���N����{�]w�n�_ F�m�]n�$��R��`��*(~Vᕼ�}�3dぞ�J�+�Ȃ�� ��N*�=�n���9:�f��q~��"�?�S�I���V:V-��/�5�����%��-�j^���,s�÷��"� ��R�4%�j[v�裏��|��W�DM�g'�t���p�KɃ� D �������*�$i+�F2�y%wQt,v����{����o�KȊW�/��bJ� ϕx4��%����Dj#�6��^"�<���#EĘ�e�����'j��v)��\�;�5�\����CM�Da�Md��Z݊댧���
eP��"IG|]�p��y�"l�U)�c[�7ҙ�������X�BQ���R	b[�����A
�)�%�4��fA:6���Ci�UO��	��|�BB�7�Rj�����
�u�%n694h}�M�6�+��F������*�qP�O�KK�3�U-�_�1S�L��>mIe[c�8v�R%����ڗ{�g(
�~*[A�YӢJy���C@��e��Q6�3l,��k��������ߓ��WS��Nŏ$�����Ҵ7�(V-1H�C��U�XWL\�4)���~�����b�m����ZX�@�����(�w��?�m�Qm��(Y�L���,��s�U�3�����a@���E��1���Çu�:>�x�0�_,����\xα���y����D=T�T�i���{�_� T�3������^n�{_4�s�Ө}���Ry0�<N;�ܪ�ّE���J㷼�-�}�z�8�[��m�6Q�{"�` ����+_�J��!�O|߃�(���/�+����R����B-�����q��m`xlM/�F�P�^��TV�ȴW��=�o�!g�D�z�*��!FK�"b����CDV��T2�Α�,�?������\�h<��x-cS[ƖV8{Z:�H�׼�5�ȧ��<�*h՗ZL�(�������s��/��3Qt��G�ÃT�f�*�Y��yHo#)r yU������/	Q��2�?@'�����d�Ax�5��0�ô�s	���	5�:���B{��G!(�6؟&ߨ������6�,��a���>=����d�����o_�p͵�U�O�tWg�q������MZr ����+?&D�i��&؃���[[W�R����B��b4<h|M~������X2�Ǌ_(���
K�"����`�\��j[������(�ָ}Cx�����k�r�=N��y b�_08Ny�~�C'|~�G��A�!Z T9��=��XX�,>$�	E��R����G���������Sjܔ��Tf��/%;�寄����!zx%!b��Jx�b?ȥT��e���-�&�`z��9���"���B�!o����G����.E1���6a�f���bbX���)���R��<Q��W%F��4O��b&���������o��
ay"E_��{,���C*�!���������X����u�[��Vر�xE�%�N+�B�o�<�?F`؉E�@�T��^
����ʁ+�䘚ë+������9dWPȂb����rDC��[c�f��I��}c�q�>o��V;z��H�n7�0��m$�ے���3x. H��o�h�IE�+���}�E�����ٶZ�"���V�%�g�D���E��_�%j\� 
���k^͇<���rQ����+�s�8�����M\vV�ǟ���ʿh��l7Ӈh'[!,!^snX_|���'�{<N�X���˲?��g���|vu�\G�F�o�zƭSA�=�xA6Fs��E���7��DSma�;�!h&r�Ց�S;p}��s�?�g[R�u��1(G�X��ͮ� �,�,�(Y�� �4��<+�((*�����18 ��,�Z %�C~�Lh��&d�3���2ɇ)?��T���(�ڷ���ۙ%���TM{��lugV���n�s)��9_Q�X'
Z�Lաk�I
���iʚm͝=ǬtQ8�j:=�����r�-��ũ�dR<ZU���X�g�u�uR"�� ~x��!�Z�#+�,Ă*ب�rK�E`��/Xo�Ḋ���U�3ް�?��O�7�����_��_�؅�����YX�4Ua|���4�-�U^$h1�Gq4)���2��1I:�!��7F�ƫX8U�"�-Q��z�m≰�����_)猻;��k�TJ����������Q|��^���M_��}�K�o\V\]�$s�`�z��>���d��
b)
��@Lo��f��O,�F�����!V��a7�/y[=g�IQ�y=�>��R�x��IֻN��#Dm�X��(.:tѪ%���7�$���XM�W�1n̂��@�?1��lC�Xǀ�[�2�+'����u��	H&���DH�?IGwG��ŴW�q�k��������I%����'��-Z�>���dՖ��N%ٔ�U��1}�6D��Ќ�5�W��U�Țc1�dl$�0<��9�Q��W�V�~݄�����L�o$j��ppO�N�?��8��҇�9�I��C��#���F�TM�Xt�z̿��=�� lKy.O�k�&C�J�<Ť�3��.�b�?�fo�K�B.�X�r�5i4@}`O���C���)���7�֢��M����ĵ���\CV�g�(�3AU��X�R^����D�阽���,E˾���S�Һb2k��ux�8�h���W�D�"P�9�43 CUOy �k�Lݷ<�ƷBA2<|����YO���VD��+#�-wf�T��==s���ٴW��Ty�[�^	*�3�E3$#�gE.M�9����D�)�llk�%!�����xeQ��E֥�s��e�Y~!Cl���6��˛%�&�/
�
����+<!k��J����\C*TI(*	�1#��S��s~?���י�&	UOR���:��"f�b=�>�\�:O�_a��G��O+���U;Ey�y&zD����n ���$��Z��K#�?U��E4n��"���_{?G4�$;��/gƛBV�����{.YR� �ښod�����7͟?��M�Ԓdf��+��H�Q���׾6\t�E�$D��r~��sP <�LEbp���z��$�'��T����b"���7��h9u@Sӟ��!�g�#��8F���Y��9%�E�,�&�4�t}�U�:MT��<:mp�����\�׽�u6>�؅n^���ã�?6�8i�։<o�5����ق�n�=������O��{�d�ƍ��w�&�T���D�&%���Lpoa1�9a���Ț���@�(!rI��	���g��_�z����R)ԉTVń�Be`�9,y.$79~�!�bƱ�:Y!���3Q�L�+��W��ն/q�����h� ����7j���˾�e�m�ehK#Q"]p�Y�O~��+��v�+���-��Z�7^�C�"k˶��1`���y�ؼ����b��C��v)U�i17�p���k� CNm�JHM,A'�'�^��c�'�������
˱ `q�|W��^��(�a����J"��K/5���������}�5�� ��7����>6�����!�EcY9�ٳf�{��'�-Ӟ�����O��v�i���\��5ض�'f[FD�F5�'!t��=R�R������ʿ��  �IDATK|<_}x��Ǫ�E����C$F[BO�ࡒ%EZc�&�΢0�^Z�|�J�m�d	��ZQ��9��0|��9F��.��2k���9v ���+̪�C߄�[{N�.�gK�-���u�p��ϸ�W}��o���GN?���]u��/]�p��(+� �k˶��v�!t���A��4)N�EL��_Oi��P%�s�,F*�����{,dB�����o�=��_,�B�������*����.�U���eL	j) <�n\S��e�b�E��G޺�0��x[K���CG<�w���������W+N:��xa�V����.�BJ8*$E]J�����x$�^���#Z8>
�(tCD1�r����%�&%E̽M%��P�6���
�����VHj,%:Q��J|q�GSi��?���jKt���el�H7�`�{/[��?��?�g����~��߽�_?;��T�����˷'[�dbЩ��j�	��LLe�'��)&�z�h�Dr��5�����)�9L�xxa���'^W��ؿ�f��F�Χ�5�����ب�=��S�s�i��q�����ZX5�5DiKs��F�E���U�|�W�n�(�s^�������>��p��܍��L�3�҇z���r���1�})
D� ̻�cҲ�FB#F���g�T�����"��p���#<�J�[����2�$�
u���CY�r�J�������dm�߱@;}���>8g!l��6������p.)�^�~_�s@	�j����}{�"�Aq�~#�c��)�(rA0��]�a}8��s�Yg��~[.��,�_����}g	ܡ�P��W�@��ZĔ+R�]�FW�.uƶƱ�PZ���:-ORM��S�ҟ�\������ ����贿��~�zvϬ[�;�[�v�(���E�\x�_������y!����3n���������Y)�XNr�Q�ziԓC���'V>�+ioU�m�(�,w~���z֞��K!�G0V�/v��C\K���?��k���J��x�a��^���:�!X���ndyRؾ�I!�祰�/L���J��gG������Gы�Mֺ�N�C��Їrg%�=lјѽd~�}������^DcQ�V
�=�P�M��>����<~�,�>G��Fk�#�2e�{ Bu��2��5����.�����6� 9�S���{^o�y�Oc��^��d��j5�h��"��ui��a`���:�+�f��"~�_�x /�1���+W�H1�>Q�)7�S�� �}ݚ����Ś���G�Ņ�,��x��\��r�0-
Z@����/�rjF�_�=�_�I��2�����A�؁x-z_:N]#]��H����s?���=#&"h,�џA���C��gh|	��חmiAW1"�)�HV�Կރ��G��M7ݔ�85o���}��;�h�^1��8���/~�w>��4�݌R�тz��o~�7�x�aq@h�0=��Y1�~D�O�q���R��)��&�,:Y>�z�]�c*���v�R�2(�B2J&2�e]�-��yJB��Q�C�аV=V˵�-�~~�P���Y�=�s`�{�+^a�y0�:�΅B4�g�������0��̈́��,jfy��q�������*�H�PD4��Aޙ@��}���c�,7VaZh�D�x�Ɍ�Y���&|}�T塘�5���C��3�<���og��G.���?��ˢ����'Ƈo�T�鞙����Wq�vu��1֎�&U��\<�rɬ�v��L�<=l��ΏG��~���&�b�b5�����6����{�"�_�I�&��5���-=����
���h��G<��o�鷃�Z������J$��B4�Z0u���4v���Tϓ.BZ=��b�ڎ?�/�k�,�d���l�"_F�����4ߢ�A{�0٩*Zp�O�Hظ�{|����[��S�q���?�㣟�������%Qyv�϶�?O� �#7��S��DO���\T�|�Ᏺ��p��h��Q���G��w�����xp��U�+�h�vw��C��Z-�,�Ks�RZ�aÆ���^��D��v*�k%���TW0^��r�|}��DI���¥~(~y���=%c=ݶ����B.�7n���v�/Nd%�Y���Z.��̍����0v ��xF_��+dO��Yq�Iy�B4iq��i�>�����@Ź,c�'�=/�S]��ո@��q���.�<��ȌS���_���~������V�`�EG�B��ʯ��OZjB�
�sd��z���'�����)��p���|�q�-#):�����̙��W��e�~����c��c)'=IG)�UX����k�w*)���&�Ox*<!�89!!W`�$�O')�<�W�zo�����!�c�9��9�~�Y�
�(ɫs�sy ���/��/_~�G?��w�m���<^��ZT��4 ���X��.��ҷ$õ?�;{�"����:�dF�g-zr�XK}�L�^cYqx�'�����1���Nr�_����h�X1�1�O,�����/|w��[��T���_�����߿��7\s��M�o�T��RXr�YU��M$}֊����2�a�714�O<?�(������q=��������o�г���Uc���]PH�k��{�`m�+$,W�IAR�bŊ�ɷ��,h%=�7�=ďC�p������V�C笐�^�|��7��y�I'���&��骫�z�%�\�!n�q���1d^h�����},_�(�䓻S�D����g��[^��x����/�QP`-�B�y0����P�ђ|���{sl�og��G����7��w�m��6�n:;��]
�zqmo����+�O) ?�䎓��i�mb,��b�԰�jõQ
�Oબ�q��5�dg�GY�x�_�����G�R��0~/#������>��Ǉzd�J���RH�ڄ��zƆ���?��?�Qu�x��Op���;��7\{������x^�c���șI�
e�=���O����ւVTƾ���-��Iw�������]-J��9}�y{���j���6Z��L�D�B���*����y�����[�����~�����-oy�O��M��^T��R����
�Qp�V���sl�뮻.�p��H{����I��W��"���o�#��څ�כ����x�O4���81���>�+���L��^#����Tq��vi��9�3�_y啗���kg<����4+U��\A�+��зU<�����pǈ�{�ޒ�I�W3Δ��h�f�;�!��� FyGq����֊�W\������n˾g��G�K�ȥ��M���OƋ��Ύ��!�Rф:T���PK�\&Kd�kr0@�!x���p�
	��Ysf��j��;n��N�O�&Չ�+tuu�[�[���w�p�	<�y��{��8P�[a�}��YR��r���a���	����7��E[s,�{���/������*q��׻��X�2�a�l�h;��*�v����z��oG����9.���줮'��kL����d��'-��������u�kf �)m�ɛ_��W\q�;���/���G~�O��d~��#'d)7��<���x|AS�2�
u�}&.5��"��Xg���)/�XY'��/���:�c�)~N��؞����}r\q�f��tW�^+�-Z��YO|wQj�$�?��u�\s�����q^����W�σ�+���(K��m(�������#$R����d��z��>
�f������M�q�^�]y�Ag���l+'�w�����y�{����\saT!�tw/����Cx�f�{{����ng�q�s�����y��Y�U1�r#�6�Y4;�fʩ�ҁ%�v�����+_�J�c���8;�.��{�0fY��9�����<�Fֲ���!ت��n�������:{������+�,����#������^�|���H!-e$��x�\&���*e�|R�I����h�<�`���8a�G��w����}n��n+�:��������ݯy�k�sϽ��q(ύ7�8��;Z�'���|��P��^\����M����m�������ۗ/����u�Y���ٽ��.�&�&s��=��me��]<��O?�l�n���mrmN?��M�������O��O�|����&"i�p���P:R���h㦈������1�&������=��1������ӎ���ۿ���+���}�����?+ޭ�{�����7���#������{��7g�x�:';��	�T��	���|�é%�QU�B�H�5I��3�C#�+_��׿+Z�+C��z��Z�kD����+��s)�����a!FY�8�c��ړa,�����>���;����x��ZI��"���7�a��o=����-�&W4�8&<�x�6Ɨ���g�]��O������{����	�w[�� o{���>���~��{�%��y�Q����dxy\v���0]���WI$CV~R*���L.8����YSa��JI�aҷysR��`F��,,g�rV
S.�=���R*ل��;R�YRuk�4�`pB��RP��;E%b�����y�m���@���x�?�;g�G�F�#��wߓO<��/�.]J�w��Y�f͉(�6'������q(��bի�#Wz���z��Fp�Xyka��%�F����x��h�sSk���^o�F�go����9ȧz�Wuu^�ˮq��R�G�X;���@�}��J�8G������m'ʽUʕ�;*b���Qf����8�x惵�����rg�(���R�RI�zŗꎇ�}����'�\J[ܛ�{T����j_<��{�������C:�8����7��(m�������W]uUwTB��гf͚Yq0΍�DԡS8�y\��%j%dcJ�n��f+��w������7�3N�2Ǥ��5Ǥ��/����&�4��1��uR��'������~v,���qL|���K�������x�~W�Egէ>���ƒ�x≏���?�hT������R��n^�#�e�m��3>*<w�7�d��g�W��H���Low<^����.���,����w	r]�d�Prz�K��^Jo���&��4����@��@�����uB3�;�Z�T��{���;z�I��ܶ�1�W�XfPƱ�~�u����gOs�1�V.��~z�;����y��ٳg/�ے���.u-;^�A5~n��{:���������k6��㸩e�|>_�h��yvM�l��`���K�=*�����54��M�D�%��&��9r<�cw .��K�,�׭wٲek�9���7�%m�?9�l˶�
m��r�i�Q�{O�d�&�(o*������k��Z�%�z׻n�nm٩����ҖqH�M�J�������[�Җ��@i+����-m���V�miK[�2����Җ��eJ[���-mi����oK[�Җ(m�ߖ���-3P�ʿ-miK[f����^��2�R    IEND�B`�PK   DU�X��MY��  �  /   images/f7330a66-6727-4ddb-8762-657115be29f9.pngtzUT]�n �`	�ww�����mp��n	Npww��apܹ���xzu��^{�쒯���P ��O�>��H�+���qm"�}��Q	���!:Hk:��#����$&���GF\�0�4ޛ`��P�~/�������B4�I`�&������n��]�9"� 6�E�|ڑ
���
Ǹl��:�$�5e�m4���>7^?�9vJ�_��a?[�BCCv�!Dٲ�"s���#�6�Ķ� �5��Q��ߙ�0�o/lF߶�&�V�PP�<lxk�ylO,����i� =�0�#�!��yU���T��gBy�zΐ�
�X�N��]�#h3�5�\�񶼷�b�l��`��� ��
���v��r�Yՠ�#���O�S�L���!�i�%f�6sB���y} >�Xǔ��C^�e̜�۹e�R[��8��bT3����4(�V���������WId�RPɒ����%�* Yr:k���H��`�A2�N_�8i��/�9��J���#dI���%.�~�bA�t��B%�/!7f���q�!(�/���Y�ǥ�"��p8=5=�*5u�ʠ�2��q�$g� �� E�Y%��2�L��8G`�$�:[Q���NP��E@(d'߂�wr��#��WDhP_ͰMܸ�B�>`b
3�WnB�_�?�3��&�����E6�N�7af�,^B�"��f�W��&w���$�F�L�[z�����YJ�;]�k� �9,A,Ta`�F�ot�i�m{_ȟј���(�?�ͅ�^˷mYa�t����b�9<:-"���G4�%h]�($D	�hoB&�������/'����3�?��ޚbI��6��;���1 D�$�r@,���r���c$~�30\���$���C��8�X�p�i��u3hK
9�;�e4�Y��)�<�����_ ���;�w4}�����2�q#�4�$j��7�՗���}�bK�}�p��}ZX���/F�fJD����Yg�g;�r)8>MȜ�B9=?48�����v�
�)��V�9��߽_����C�׫� ��e���Nû]���K�S�i�D.��9�߹w.D��3�1�u�,�GS6I�6�ڪ�1��z���2+?d.X)�+�'S�	N��M�"��ú�_)+?��w���IEP�5`���-zM�BQ��jl�#�Hf�\!�|}ڲ�:�藀%]�D¯@M�(��i!Ĺ��U���:�:���U���L����Q����XI���ղ�����s��!���Z�9��wܷ�[\tTu
&>\�W0���,��QP��s��L���^�;"y�3����O8�3��������j;o&7��jw�R8M��%�d2���F
]�Oe&n� ګ��C��]&ڐ���&�NrCg�`}Xy�X�&��#��9�/��j�Rc�v1�����!�?/���ک�����͖��^g���~ѣ���~hm��^/��t'Z<i�ef�y�ˊ%�����)�dlK��)F���d:��q)�?�'ݿ\�\�Gon�dba0�$wyݢzW�{(��G4��d(���=d�'��ɜBcebB���Yju���LY��s�4ڮ���N
3O�2�ے��w�Fܟg����J�¸�I�4o��H�+��u���9_5M��`�L+�j���7�"`�������w��蓻�lT��iJ��h��Q�vaP/,9Α�Dq�:���YI�v��ƨۭ��;/X�+�}^|�c�9��L\c}�;c6�hh�^O�Y=�Lh�G��Hx���a)�����{p���:6Kݏ�/���5���e�Vc7��|;ܸ{��k�ϞN���7iA�!+�[I�؍�o0�Ũ�ϖ����4^�\45 �cS	�@�F��uf��>Ve��j��D�Z�>h���r��:����&����/ʍ����8���g��۞���3\5��u'<�aG��r��5�IV���(�Q{�+\<M���ׯ_-ll���^!�Xr�/�רk��9�O�_�S�#R�˿:������n���EY����4)|��K���i��bs����6�|�y��5�m�x6���÷ۏu�J5O���_?�J`5dƨ/��1�D�ғ��|�#R4<��E�~�F�LJ�P�����B�}ك}��.�K,Q��	P.�|9v|>k�M
���NrEڶ?mq�1o��m�=/��s�i}q�Ѕ�?����!\�(�Ps
�@�iQ:4IP�������Z�-
���XkAX�k�|�K��Y��o�je��ݿ�g��
gꈾ�}o�����23�����zf�IqJ��/��ֿ��B���z8o0M���oV^i�G�6�"!I�S���g����P��#����hr�����Ϻ���ꂏ�yD���p|cf�˹�s�P(w���!�c]&o!yB���.�}�w��E���F�|^e+�-g2½���c����
Q9�rx�ta4r^�}��� �m�Ԕ������P<y����P|�-''�)���z�K���|��'��6��,9��p�X�wS�UgkZ}����^A��RW�����Ѯ���*�ܞ;�:�0�A6�P���6_/w"�N���ҍ�2}��W��yyw�x����8-���鯚1�È6+sPY%���/x�ץZ��Oz��q#�!0N!�F5�F��_�Q��Q��(�8J��q-4mH�	Sl�;9��X�D�j�5�c-d�䵷g�� !������98���G���bOSш��01��9�=@�[Go��\���@���1eKQ�����i����{ �'��7ѽ��_tb����+��y��iI��Y8����ţ�uژ	h�@�[�aD�	0Zc�r�f�m��a)�x&Ӱ��gt��P[( ���˙��É��D=�A:�h�����K��u�,���Ӻ���u_yzz��mB����lQ���|�+`���5{����TLP[' -[w���ޭ8t$&_sɕ��Π�_�]�gQ����͹܀��C<��F����J�B��c�*����c�?����b3BC�zRنʦ9�{u�\���Z�V�+x��a��+dDf��ᕨn6|;�J{,8=f8,r�4Et֕��;ܽ���Rę�C:8�-b,�8Wf�Ջ��$#�&s��v-�9�R��	 Kw����j�>̔�S,�,5�6{(�P�(�\�Xz��GL��@�?��Zk�7�<4<l�:��������������T����h��1&�|�EWwx<�*���1}w�N}�������m����
y
�����ު�ΰڪ�Ӹ�PU��h
SRv�(�}�N83A�]"���J�誛����i���b�����zzz:����^�~h�#�>�6�P�G���)*��J7f�O�����Q���>8V�|�:�h#���m#�ئ�����Q�l���Jcc;�)g��G\��E���͏�Z�z҈�潶�b{�p�0��W� �<�'������dE6�oq>����/�TH���FN]��R�X$�����&8�	k�[���;[�8���K��~hcͦ�0cy7GhN}�,Z���j��8�ٷ�����㐴�.h/�B��L�]��%(:���_r��1�񀗗*��0��S=���z�]�7�0��İ5翤Z\Z/lI&��{0��#LFZ;�#J֦�V�Y-�Jv�55Gb�3����n�>�϶v�g65��
�J( �ê��	��XO�Ozj�^�klLA|���:�^�� �b��ϑO������>��v� j��q�?�n�"��e���X�8��0�/��V˱��� �Hg�����^q/��ڃ!��� ������[�Ewb{A_�aGd�p�J̑�2?T!�w� I�+�nB-))��>39�g������a��ni�2]�k!���$א�P�8�F�Q/u��N[K��X�=�hd�ܤ=��������e���D�o�.�.\	�{�L7$fjT�%��Bُ�M-��JrT����j�/(��4W��M�U�sD|�o��8�n\i2�F&����3�ug5b��̲�;#1�~��=W�a�;;���T���cu��3��S�d�܀�6Å}�I�x���м.Kh��:�6.
�N��>�#!<�u\Hbd�ٙ٢�𣅄����`M�'}غnޟkd:ct[8l�Fc��q�^tc��Ew.����ģ������k��t�Ce5F�d��y|T~~����B����CN{Y�h�1�P�2�+z,��	L1~�>zR�����;��3u:��7��/�eU�5�s�c��FK�e����ǒ"�ݍ�[��f��H�}��jC��[-�^�T�d��j�}���*�b��2�k-�����-zs��R,1w>�Y_U�ͤ��d�4��ܔ�f-J4�B]KW�����Ա6f��>���ze�<��������aK�d��l�㊶Ɍa�{s6Y͹�]&�$���2O��P��}5L--��I����>�-��n޻�IR��=�h��][�����d�����b�h5�԰���|4mgm%G�Vh��C%�MЃ�x�J�	P�#f�Xy����4�B��Ҏ��RU�P�����~���YK����k�e0�M��A��yq`ۯ����3\��]�v��ҦqX�����Y,���D�OdB�9��9V~
��DC�J�~͠��Nf�Hň�E:��[��b<�[�L�I��B+��S�%I�S�]ed(��c��+V`D䖏N��$퍦�w���$2�͊��5~ŪϮ-@����i�T��@��`<�X�s$dGX�KY2hh���&X��~`�m�NV��Ez;`��T����D(B��|��� Wf,V��}Ã���m�8�JĠ��O_c��ʄ�^�8	=g�%���jw�xB���o�J>(���(��O��ϝu��Y���a�w���7M�L����}�c���B�q�E�VM5x��BCq<�5s8L}�
M�_$�t�MW����Ĳ#��s�$�-̴U�����H���?��Qh�lU!Ę�t)x/+;.~�6N��������<��D��CyEAI`L %t��Y���	}>��zh�zPep�{�ab��U��������0���D�����y7K�<��/&s�f�6�"S]뒅9�h-{�sޞ���,a?!��c������M�6��@��˻ �m�x2�N��c寽�n!Y�t)A�d�rUb���29p�'LZ�o�b�$�.�gn�1Sq:����U���vi�Cҫ�WlB��8J��%�o_ $~T�v�VV:ꪈ�E�AU��^����P�C"4���k���R4��7�(�lk+0-�� OT���Bo"�! ��bt��v�����'���^����R�ܨ8�f�V��w�>�_�WоN#�����8�ڗ>�!ak�b��Gjė��1��	�B~�}��mc���҈;�bG�3/��tT�؇�mps8Mu���{�hһ��}���m���~~�	��I����h�tT����MP�d��n��E��!t˟ޚW� �o��^�Dۨ�6sLtH|>��'���]�=�-,�����`�"���^�F.(��HR�<�#�ԉ^�=E�A� !�q�Z��WML�X��I]r�$C���d:�l�c	��g�|[�:�`$�Y4Һ!H��/2155���7b�PfV=r�t�FI��_���0Mú�O�Z��T�*D���S,S�n%f��ߕ�N�!S,Q�fԖaV	1���i�~��,�2}:O�^��<J�J_� ͒��#t`W�g6�t��X���a]��+2O�$yN���5П��$R�#
qLe�R��;��X�|����R3R�qJ���z��ʐ߿O���d:8�/�������������n�>3�U��l���/V�����>�����;]s�dA�d\�;��^MY���?7O�b�������o�B}NLSS,��>-�p�/������_<��
������+V�#�R.��-D�p���E�C q�ŧV�������b=���Äew`艚�M�����8�^\�����J=�>��%	HP|3��`��u��#82n���}�1�f�;ň� _�S��/�p�;�m�NM[�AZ7���Q�S��޷C��f�Jô�!�x.�����U?�v ����+	���\^E;�_���gӎ7<�"{� R�b�u���E���P>VEY3��kb��o*U��)������ԣ��=z�L�F��8��z��8��}K�G__Q�rշ�~.�	�*fegP�w���*�	�G���F�?������ �U���
8�?�i����Ã��2���')᳸�����nK2w��5��MŃ�+��e���Q�����4�j��*�����t~�B��ة��OE��ӥ���a��bG��Ee�I��v2������эG.|��k���q1#��%l�	�z]�^/��x�q�D_�p�'��C���'�t[�=_��OH1T��{�f���6���_ 	�W�t/�+lj�E�b�)�O�M�U��R�'q��b�ը_{��>��dY,P�!�o�I�4�U��{!��N�
��!�o�bt��n�p�D}���zf�Cj�����28`�e�ZW��j�Ӧ"z�ޱɶp!��%��ސ��R[U��RU޵���#�7\�p���_�u������M��a)cp�ɶ�	={���I������;1�T�#:�}CY�3�8���DL6���ѵ���8��۟ZʢЋ�զ����1~Z�\��#�X�ٽ�!��=2�������S|������͓��V�-���o!��Vi�YW�h"&.��A��'8�%r�.Z(�'�����;��I�:F5�gJC�l?��Y�:���~�V8�U)*�d�a�m6���lO(�����:.ݐ��aք*����Q�	v�e����J}�sm�3�\�L(&�D�+��kR���W�Vd��6���P��N�IR��nr-j�e
��6L�W��zU�����x��,ި���f��r:�-n[q�׮Y����|q-�
��Bl�2${]�X�I����+����i�3�9�W�����L�7-��6	�ǡ���A�0/����y���5�����u��ɓhFH��S�I$���S�j����2�"��K|��z!��������	����o~���9-d_#�k��*�?��$J�S�.:<����q��{Ӻ)��E��������J�݋?�-�|K�UpY�����>S�r:��Zd�}%A��	/�g.�O�O3w��(T������e����:�:��w-�4����W�tÇi ��Bc2dJ����K��I-;j<^�.�f�qr���1���|�.�:V+�����+a������B������ �Sñ��~;YSDa��_pÝ:1Eoث1&|��o$�p�%�_l�&Jv�庠�X_��!]O�܎?# G��mԜ��&F���R@Q
ho%�*qCMys��s�$�Š��f�_�l���6spk	�`���Г{�zt�0ѩ�[���,:�W'lAuw���<ҝ�1<_I��(��z�
�)�2�����9B|�,s����ߏ|��6��x�r=5�h�N��;�!��d=1�fuZ��Хj�\G2��:��ܼT����(?b˳�5�KT�J�\.��)j0s�LY�+)�;���z�,O���Y�[")5�f�ˁˉM
���"tGY�˩t�	n����|�Ҷ��*Uh�D\�rwmq��fc��/s���2���x�T1l���Lh��& $d���ȥ0[�'��:~5J"�����������QaB�����Lc�{�QN���S�͝�G��4�cؖܚ��:M��4A���_:0ѯ�������xlq���0��7��K�_�S0��/��G�a�����Q]6�bEd<������s�~ZM���.���}2�j<�拵���LP]��\���7�!rt�tWy;,#9'ᗗ�����)Df��,�@�7J�d����IVwy��׎����~م��ɛ:���%�ŝ����Zoo�޲\���*C,S���-�R+��S�Mx8B���4VlYp�]R	e����6y���	�㛘v���h�$���Q��Yd|Tx_� 4tCv�\����3(S�c���>z��ٰ�+����`��h鱦�#�o��'��ͪ����6b�Yv��7��'��>Nd�Zy�7�w��a�쮃Vp/���.��i��uə~ �u���ۧ?�V����Ǹ�Qhw'�t�ǆ��f�(G�'����h��ʏ�I�=(ēcq�؈��w%ae�0T�J@�]O��V���ڒl~����S���(�Fv�lf>���_F�l���n-l��f"1��|~2Xs�}�B���B�n�xHٿ�H8
�{�rs�j�����o0=�8�{y�����$��k��hUO=b�M����H�C���#�[N0�&�y��+K'������I��Y���5Ob��
�jb�oQ�`A}�-�9������
i�|R,Gg���PK%�:��oLqж���_��a��~$[� �?5��I��GR-	^�oٖ�\Q����{�|�t��jv�ONHt�m]��T�u-��(^�l~�����U0G�5OK/lE��o�KD�$�����
�w�������]�8��
�Ķ����ҝ���&V�$,[@��E�=�Vi|��m9�T�����9�U	�8����s~�G$�d6�Ͱ�[���֬��c��������P�k��v"����j�>�f�$���ĝ7�1�7��y��N4�_��T 6�ϑ�V������q$Rb�?&g�Nr�ˍ�����2�l�aA^�;�C%8�WH�S�,� ���f{�h���ׇ�-�|�@�e�U�5Cjn6����0'cwd�lp&��|,���8����mS!������L��x]�boHi&�mp ^�v�M��/�t�nc��!��4�1bS�u���P�ٲ��"�1z	���Mz�z|De�نv���sb�<y���Zw2���j��-�+hՕ�la%�5����/N:�sL�I�\.�2����ދ�^�������;8��,�y��h�e3����S �WC#�V�`n[nV�_���Q#��> ��1jݥ1�^����q���pD2���	o&�1U����-N����������u0�nɂ���U�0{T�Ki����u6Z;���j�n������<��/$���j�q���W+���}��'��K����x8��ӈ��\ʊ}y5�]<�cȤ1��.D=
�0u!|J3�E�x0�)o8��dؤ6`�h3Y�4\��'Xg�9����Ei��ݺ�:�4����!Snc�n�ܯ��ȋ'�4C±��8���o m7�%�_��$��&�݈�*�ѵg�)����k~��J��^9�<�~͈$�m�+����/�Fؾ�}tYWr��؈���d�Ս�fb�\Cg��Aתp��*W�~'*��d��
�D!^��=���;!Ɋp�ޮ��������7�gv�K;br�>��j���P"�,�.-��*�#fq �N�ĪK�O%+9­��h|��6��r�iߘ2�lZ����$���va�|���8�~a��c�)54[d�s����GJ�̫\�!H(8R٦N��8	�"�v�L�=;�h�D��j~:�دT1�H�#F��~�:d�S�bS��_�����}�^�=q�p�~��y���맼߉�B�����W�Vx��������{XoD�']Ha�����Lk�ԭ!���gj�4����4��P�P������2���f���t�|e�] ������e�P���X���g��Uh#k�@��)���v<@Α#'E)QW�n����<+s�F[h�S!+���lί�û�=��^#_���z�!yS�,A�����?{��Ȉr��lv�;�$�D� L`��ߝ)�As�Ț�Xr��@��T+FW����Y>?�쁆���A�!5b �����'=D���왣s+U��QgE��������$�4&�e-�r������c��Ի\��^��\O��c�o� [��*�yD͝�oe�6�p�N���n5���ʟ���s��q���*#����n�&�ژ�'�p)�=��,ss<�p�<<K�����=��4tak����Cr���������eӲ5G��E$��P��)r��Sņ����ZV�>�[?�ݜ�1�W�2P� ���G����O��w�27�K(�Ǳ��2*jכo<�1W,��9��g�ѩ�c�/��?�2ㇳ���+D��o:�KG�3q#�����ژ���EEl�E"	^KQ��^h�AB!��1���̗�������<�rA�U�G�q���W�6s������:�KL����<���u�io\z3�o�l��i��InM1o��\��alX��MNF��8Qщ��e:����3oDp��#���M(2���e.�L^=���0�b^�Z�H�w�� ����WyɎ�ty���q��uy���l���O>"��{��F˙��S�]��D���\�����R�����m�L(��ct�>< �6CϹ^!%n؅i�X���X�J���wC�,���VV6��x&=z�(�Y�(b�!W�B��"�͙��qmF��0)p�����������yS��.S|�j�5�2M��^Y���ew:b��Mо܌�8��" �\��Н�؃���O5Z��7�oa�ۨ ��S�X�_00�^���3���O��<�74jZ!?�r>^�i�[|U��	'����=}��K/r���-q� qp!��xJ�q�QMi����V?�r��~E�s��m��%�<F}�q�4�!��2�u��4��-�\Y�ndw� �٩)�hn|����7�F�������g4�o�w|6��(�����B���`g�"�@s�J�:�_��A�z��F�	�Q�M4��9�a�O�2�q<@h����X'Ż�|w3����1�Q�!��{7GiP,Il�/n�ٸ��zJ:����LA�!4�C�E��p�H-:1u��h�֝�oL��hMgϺ��;�	-Wu��%��/����V���e����	�կ��<A����t9��#u�kl�'0e.oY8J[�m|oooc�W;��l֭��w�]oX]ﾣ��ff*�l?&<2��^��f)Q *�'�)'�|ct��`3���U-�����ɓ.�9�����5�|VQ�sУ^��w�R����v���9�%q��!É��=�#QQ��uԅ�����}h�^w6\����D�j�U���q}�������D�o=!��cD僻(��@���B���
���xz�0?�~P$�$y:%�y]t�5�9�J��g�����^`顮�o�PZYZ��#Y��Xp�M8�#ލHG���s�c��_4��Cs�q� /��b��ř��Lb"���lAw���SY�5E°���[���P�Ũ�C%i����-/G.̑��MAj>�@����4�{�Ѐ��!�
���]�:W����Y-j͉�))"^���/�yfC�.�PF�O� ��3?�1>���x^���q/5]x��l[�!��[~ѱٟ[LX�D˗w5����-e�cd��1�(
e��\�4ݙ6�#R����u5L�<���L���O]u��9�:��.³^��#;0�(F__?���
�l'����Ob�1�ЕOM6�ǥ��y� ����U����ҁ+�Y��G7��O�)m����sQRHeE��_�^D��z�n���ck�&Z�P��db��Dp�KRf�.�;@��K#��S}���{�w���tT�����!�.=jTƽo�c��+��5�x�7(��/߫���b�\L�>���"�a���A'\]9�k<�RC�|�a�o�X3�ybj�ѷQ9R���;�z&�'�߳����9=��4��Tk7L��P��G�v��o�C��E7N���a���C������ל�қ�g	�!���jZ��gIY\b�/o��<���WO��p��N=F.f�H:,�-y�2+�&}��J0>�'E@v�>!~����I~f�x|�k�E�@�R9�Ӣ%�|g� OX,b#�	P�9������m���̺p�t�R��"-V1�Xy@NE�kNv%��?����=�ͽ"����xv;	St���Z{�Џ��"u�GZ����LeS�YG�֠@wꇪ�d6x��=7�hb�Fgc"�����D$;���l=�G�_��_��;�'�o����v*��TQ��B:T�g����|�����?c�yT�żo���d�.wb3�Y����_r�%�3�X�d���ψC�xQ��?�AE$�3.A����Q˖�J"2~Fڮ�V�
��CJZ�����y��,>�\�>��Ul���*Zl�2I��[N��m�͆�Z,?�����Rhb�����|��g�#{}��eR��{�HA�����d����*�-с>�|#�#艿�E
'
��ɔ�^Y�R��o�?�Z������ ⡄����	}����M����5?���[��*��ąK
@��N�Ekj놎]K9����-��}_>�m����7��ן���mԜd���>f����f�K��q������0��I�oVg��1(B�f���B�|I+���^�_?���6����G�6��}���o��")C�e_Ry ^�~A���޷��N�BK`XN��T$1-į?M�N5,Vd0rC�M��X�To�����p[2@��8v"�ڣٛ�m�C%�s�M��T# $ە�z��j���@��EmM]6��\�h��� �oG!	L��4_m����8��ɳ;�}�я�ő�O's"��}� ���e�'��&@�t�	k%�FĀ	yj�R�8sǢ�׵�gF��8n�;X�̢�o��8:k��bY���-'�4ǝ���[�_�x���tar���*T!EE��k�V9��
��̬�1��qC�K�؈��wae�%9����H	�_��ﰤҥa�a��;���KX?.r�Jj�T�:6n�"$t���5�����w�GP��dha �PfSq�t
��U$�����r�"�4��kq��HG����Y�;�Z`�4�N����
T/�E1Qk�2�#��]8M��C�:1H��]ԟ�*����E�H,��On�f��M|6����]4g��^gɚoQ+���#�<�Q��=�E�׾g�n>���_[�)�
%Ao��Ur�&^�_��_/"4�Sp`�a��huQ�`���`�S)܌��l������w}��
�V��p�|�Q���$"�<�O��]���s�`�ۂ�8��jP�'����k� ���.|)]]_Wc��	�/��.!Vǉ�q�{Xޣe�7�W�Ǯ�K���ž����?>Y|��ph�Y�p`G��B��C�^w���׏x关x��z'�P{yQQ�^F/SR���n!�e\�vʡ��⽂w7-��`&\�G��)��Z[?�Ƭ��<=Y��_��6���>�kJ�X�Ǽ]��t��7;�u��EZ���鞇�y�˞����|�-;�'�f���4�	ޜg��K��v	i�k���^�W4uЊ�)	f�y���="BTwz��?
��N+�q\ڦ���m�!I��A���:��ڝ�T�.^�a�t��XBn��\u���u߫���rv�ߦP�5�_�6Q0X\��7*�_~z��[sy�.�ZiC����-�>� _������%���ӎ����� p�"����-+��p=[������e�}[0//�|U}7`eE��$@��=�a��wR�[������As�{��{7ɔݕ4��yT��<�#�j����������5�u�t�O��J^���C�
f��$F��0�V�M�L�l�O���lӶTS�
��������ǛS��{��qꚻ�6�0�3ڢ��N����F�@:���ZH��ԷG8~�n��A�!3V�M�J�%06rm����ƚ��D��B�v��I�=dPp1s%$�d���ޮG�%wֱ��x>�6�?A��A���[�z]O�T�ǼN�1U]ތK��cR;ߒ�؅��D���\;��_,���r�,���x�٭�hj�)��K���^������n��ү��G��`g��i��z�&6��b�0�9���_(D˴�i띡�{l��5�6�r��kl)+�u9Xؾ��Zj���v֟�8,�R?p˒5l�2v�F����Q�߻�N�˰E��O��DR���ĠU�@�^�G*���d��҉�>6�(g%�!ApP4����xzVQ(�ᗄ�4(8�F<8�3�S��(|Qȼ��"��%�z����V[���B#Yډ }Z����Y�u�^D�ڈHU���P�RA��ǯvK��>�.��@�?�}/�5\m����A�Sgkv1�m���>P�R7�K�� ݄���;:^�Ŗa'vQ%�6^��=��R0�|�V�P&_U��������%�D"Gb����b�%��Y��}�.o���k�U�����Od�ȦAv�)��×�4���2�v|�̵�t�uI��gq�+D�:`�� Q�z)-��j���-�GiP��WNY�
��1�.Y�:n&=̎�]?ߩ��������`�j���V�<_tŞ�65�d�3mx�W8�G%d�
�՗������o�2�b��i���K��Z���m��^�������E�{�6b���E�Ƕ��{�����5�X�u�����i��T�jkkY<�L���d�����a�A v(jѫ>4�����a���;`ei�;_M��V}i��Î/�Q�.���2Q^l�H�Ã�����u���AO<����ݍ`�1�~6H��{���l����3�K�9|��̤M-��q�1�CB.c��������N�S��
A�.}�|�s�(��k&L��J� m	�Lg��]��ep��>��OQ
�=0��٨�d� �No��A
u$%��߸0ՠq�PB��x;*vv�[�F��^�?���4��?�@)�F)�b����G�����'���p (����,`�c�����1�Ր����כ�*���A���nn{ㄺ�A��[=�>K�7���D}�tx8B�csI�;���%s�8d�J� 1	��F��~�x�,�����Е��C��������kA��0'V��ts�.Q��
9�z�eźJkfK���.�hyby�}�m>;��y>�g1T���+ag[�K�'�����Z��g/�����qwoW.��0�-���(8'g��n7Q�v r���=���FK�q�i]BbM�r ��p�\�V���).�k��-�Z҄ZKҦ�/l-j��Ŋ���~��Β��o�`!$���8�j�W#����\�1��A[Ԭ���""* �l�ǩ���in֜�Z����|�F�p�ƋI�u4l{1K��p�(P)���kS��{���f����Rw�dJ`�Ύ껵?�Dq\�
�T;#V�s� �8m~�"�p��@��y�&�+d*�}EI��i�J�v�����sRZ�3ϳ�*����+A�2�tX�<��% 5I�c��]��J\F����q���jd�/)W������I�։J(Zpշ��}o��V��d+F6��ep��K� Q�qς}'��ϾN��	5��,[7����#�q)s5K;;��&\�5=�n�7^_w��
�s�W��b�Ji�%�u�����vLQk{���+_�k?�q�= �&#�4&��+����C����.ˏ�@Y��U��#��z���(��|�6#Bݗ�����Z��rS�JHȬr�~��������6�T�z�&�zi��;ޖQ�d�g�O�[Pn�|x�����'�0����xx�3�auK\��rQUhd���ճÞ0�`]�hС+�d-��L��ǆ���`�F�v�V�I6��N{�+|�֮���U���U����z�2#�)��魊$��d]UygfQ��FYLwZq"�����ׁl�D�K�H��d�-+��ѝ��|�:���5VŇ��PS���y����`_�r�y�k��BT�F�gk�}���ԆF4�(NM8Gi��}X����Ub�9��H�?9B�n�������rb�/p�d�� t�ϲ���,��GJ�#Ӌ4�m+&nL.ˤ�*R�ë��_ya�_p7r���n8)|E|�p�,��5���(��z�)���uXvL}{����/�����[����暛r�*�5_���_�"���n�KS�;��K�}o0����Q�����vO�1e����n蕋�+���8�hK)�	������uU�	uh�`jތ�m�R�r�a+1������Wb�>�ٚ$��Wj�3�PFGZQ��.���d�2yy��M�c����d�DZ��{ˠ8��[4��www�w� ��!�w�����@plpww���έs�Nչ?�jj����ٽ{�^=5��:�\�3w޷�ܓu��!���<�[�x ��]g�@��=W�A��3h���đE3bY��`���_���ßŅ�ʕ��=��puO_��H���K�G�=IB|g%�L�A{>[[ ��'{��^���v���)�~�b���:y�]�b�'�BGh�f����~�ȫ�Af� �=�����a�����>j��)�{���sk�1y1�dh��G�Y^%
q���2�<-J�[�,���7�Y���
�D���+C���)����� }�"2믄Ml����Iis=�Q��݃�6P�]��2��!��S�@���u���qa\w�0K�B� j��P�C���[=B���6��R����fˁ��ܤ�_Uc��C�!�tJ�}T�a���T3B�����@�~�*l���@��ȃ��?� �rl�Efa�;��@h�06���oD���I�~���h�y����xZb�o��br=���wP�8aNA��
���ƧkY���
B��t�JV�����Va�+:ɘ<��
��5�x���~�C�h�z�X	A��n�cT:�C�8�<�b��l�mj�~[7Y`?܆JɤG�:�"�4Z镻����N_`e�K)�k�j:�p��,�.���~���(�71�3C�K���oa��}���K��Z�J�W�)ṝ��1׾��)2�ChSLE���'�������F��K3j�7`�C��/f�"
�~�������������c�nL�Hʴ��~�><���J-w�I*F^䰹��k�2�Ij(Y�K8���X��s�U����$�W��6�!-������=-?ɘA�Q��8)�����_�����$%��qv?��p�S�~�F���xl��0�~T�jY4��D���rx�X���E�	����	�-�/�	�����9(�R!@��V-�y��NgkMÜK��Y��Q
���k���	(��\:KVj?���}�,V���,UZ[�(����!ZY2�s��O���i�~�&х|1�y+���
t���suI�s��ެ>�F��.@�+���{�S2!�7�� d�;/ւ�*� vy��g1B�}5 Չ2�e`ט6���K-����6g��
Yt��9��Vh��b��Dyݿ<���2�/���Jz;Ylpl�C�;�����}B0m��)�[��Q[�ܶ1�k&����Φ�f`�pBȴ�I�Y��c�(;��J�6��g&��Xo�Z!��$A�c�d��x�h�my��6��W�[���,�>e��t?���_~���J��Cp�%���[�����2R6:��y�S��\u�o����������~4���*v���UM���G�V�v8�����k�u�oc'w��_u�_��xH����Uڼ���4�#�v{3���U�r��V��T�r�ž���B�	�T�nA�]�|w���d���M��+z�XP6µ�JP�7�Y����]p��Bx���-'w0�6�=��w/pcP��Bf;u���gZL�u�-�[[[,�0N`�_�Łd[ΰ��$�0W3}q2:��!zXS�}m��<�Ň�d
��!��qi�q�NPdd;��p�=$#�96\��y�����C4L#"bbѣ�0��:\J�$�I+Z<��� aoM����s�Nm2}����׸�܅�C�� :���E���0a�'��,=�H�-���� J�A��?}�D_�-�RR$�O�q��2���t�:�;�Nb|i#�hVw�lݧ�^3�xYjH��x���ᯮ����Ö'������Ó+����-~I2���m��'�a�*�ha�
=<��O2*)���1H���6�ځʖ[��)D��Vva+��π8�3ǿIv��D����w�c�f,�~⢻�N���v�P�ys�b�=��(��nd�	��/����y�'�b<͋:0�`�P�W2&;�s_j�C��v3H�z;��j3���B�����&$�r����p�t#�V�\���,���U�ɤ�Z��@T1ߘԣ��_��r�#U �� |4�y@��ޢ�v���Z��w���0�{�d��v��x1Fx|�ӷ.�d"}���'�4v#T/"��L�9j<�ҁ@L��3�P��ѹ�ڊ΂<V�|;2<�0��]Ќ3�U�6U_��⫱����1|8@YS&ZBS���K��	���bhce 6��W[�������%�?=�e;W�\9J��x����h�G𑸞,�B�1ݬ�q�����96�����֙-~��IG�r8�����|����s�؛y�ޘ���k�JT�q���3	�t�2����g1�OD尠왦Ƨ���fƂ�=�����*vB��k�a�n�S�=g��N8ב|='0���vW]x�xY��ãP'�4U�g��8i�³���qA��tH��{�8�D��u�Ʉ�^2�q�����D����1�4�r�Ւ���J���mեΔe8N�S`�=����M�"�<��E��S���B������Nw����G)�AB�*߇�'/4�ᠼHd�N7}m��d�R��t�W�St�8tn�A�A�n��<�d�5D�8�޿&���6���ORe���͓�c�jzJ���F.-�;��|��k�_�Wi�i8E�������S�3��sR�I��:�Z�P�oQn���Zw��#d�;����e����7},�2��\����e��G���Ŝ���;d`ϝ���Tӿ!/Z�z������汛�I�VE�s��'VYc?ԧ��B��M�ڸ�|X��8{�)�����<P�Ѧ r<���p|\�?v��u��/>�rL�\�g&�?r�bį�/�ۄoU�������y�ⷞe��ӗ��^����"��7�-p������-vP���=�K�\e�g�|;��K�D*�I�C]�K)cߦ8jR!��v����fĸʔ������*kv	��K�N�p��*� %�ל1/�rC�4��y�t�oc;�5 �u[R��M�ZQ��R-~�}�_3���<�^�>Y_1Ru�[�����f��Үh���}��h@��'�o�>���:���ŁC�8�)�>1��38 [���wph-S���;~@�C2ʥ����Ć�V�$�% 
J���"^��o�ϣX6<��!��R[�L�_�`��{Ha��.�g#e��㙬�y���_������ ����Ň@g+ct����x��Op��+D��+�imm-?>�R�6N�pw�G6y�e�e�:�s2��D�r� +	No�2u
�>TPru}on�`J�ĸ�-J�6�H�)Rf�F�'�����ޱU���q��9T�s�h*�H�!�����P8F���o����:cԇV%�8ح��X�]�c�v�:���h2�K9rݜ�+V�U�2j2�k�� �4 �������y9���ȴc����p�,vu\������!�}��Z��G�-���`�*�{<�ݐ�|��!U�����R�Ks�Г�n��䈹(��nw�'�����>�E73J4��������b/O	�-�Ǽ�i���A����]x��D�E	-�[��j�G4�z��U��P=1�����(ci�y"��V;EB�v7!T��&Z Ճt��aa1,q�}O^���~�����͚:��J54�.S��s&g-�.ܑ^�f��sk�d�!Ϙā�~�Cu��qr+�3�Ӵ�I@w��1n�1��aj���ۡ���.��X����]�M�d��������Y[�P�87[���X�z��t�p����{M��YH)�� K���R�-Y�q��ծ�'eZT���)��@��� 3(���ib�'{z��}(���*c ��`�;d����;s�~MW��G�F�������
���`q�+C:g��[���Q��ﷅ7ї�~]F4��[���#�����T1�zi�:��O���=.{Y䈸�C.�8W�TBp�qC���MMܒ�����X�`Q��*tT������d����� U��N��#��;5�)�Ӷ���?5�[5>�+RS{p���LK��_,�z�d0��9����T��u�˝��a��?���ml�)��*�6���uyJ3��!�Qwq��afW�����Y? 4Qw4�2�&^�G�#k�c�ʟYd�����9C�h:Hu�I�uc���bq�u��襬DO4H��rE�'�d�l����#�,Օ�V�l�9CjU~��ulů3�d5ND��0(�2�-����V�l�w<𸸳�B17]Hr�:4[4�W�ǈ"��rx�{ /ö��:ڬ$�a���?6)�0;��gY��x�����A�o�$�gd���{���Qnq{C���Z�on�Ƴ-^�;D�FE�^GG+���E}L�C&�y��=�`�E��$���#��G�xr~����QG�ۋ���AC�����dy���}�X���+���<���%�����
Sǯz��f��'�7@!d��7D\��ܚ����Ħ["���|��5[JA^R��-��2���]:/�Ҏ~!� �2��p���I����D=uc.?��pR�W�y�1���|�O�*M��|�u�v	f`%dG���\t���	B��,������|di�5jzM�~|��cí�I���n����
H�s[������g�xwk�W�ki��~���+83&�����e��
������[(?�_-Q�(�p|˓����$^�<��Q��~}{���͗�xd�Ȕ�΁=�z��'�����\{r�i0�Ra� 0�����q�p؅!��~�L��n�Ϳ�1aWw�852yzz����A�S.L,���O��,�hy�`�t^����!���m��®Y�W���Wfx<1Q�#�xOh��I��+��p��鶌�Z���n��/j��('k�����У_=kSK���[��nO6�1�TD3X����B\��c����.P%]5�.+ёt+ѴTW+%5(���K������x�i�d�ZWt4vKP@��q���׆�e�wg��Ch���)�|
�������5g�5s�wS�c~i��Պ%2`gd���LD��`����Z��LM�����}v�.C�\����]���iIr7��s�'���j������^��b�j�ٯ�w��ٙi��sU�H��d�p><8�TǴ����|S�EE�xx{��h��J��w���y��g�M��}�'��p�����<�#G�<G����v�o�>Y.z*S�bJ�S���-�7�W�UcDP�(.8��L������"����R����fMR#]��JQ�p�!�]�։忪���.��x@��}�-��1�o��Ʈ���%ZK��Nj�+ᩛ	���8��@�*f�����as�p�%����Z���U��o*#l��������FH�q2�֩i����?6��Iqfj;�M��^��к����DJ��F�͛rs���*S�ۦ����h�4���_H��L/�����Ӣ�_��	;-�E|� cw�̤��������%C���Ɵ�w��M��R��J.����oK.�[�X��FS�P�z|%=I������Y���\�_;���L�%!�q_�����8Х�U��`�����l8f\N:r` L�V�o|���V�>B�S�X�UF٘���#A�l�嘞���:��ȋ>/\|��̙_a�JQ��SW
��D��)�Yr���m P��@���P��|��T�y��t)QCsB
��<?�CC p���A���-�W9��r2���+Y�=�SAXl:���R�����ab|�(�x�2�HVǓ��[�b�;F�r��NV��Ί��`�8�8��_���i�`|1\�I��F��K�׌�ٸe�EnK�����m�a@�v3������W�c<�Q�l��vH�R�@yx�AWwn�{EV�\�y�(:�?#HAK1��|3�+6*���Í��b� �Ǩ������&n��u����b�`��;�w97�|m���4O8�~���f��9m��\��?�*����[��m�\���[�T��m��x!���g�&13,��Cg�v�����⸌�KAZs�0���9 (Ef�[b��]��Ӎ�ș�5Z�]��|	ݰ|	�2j���ny��9�/p�ἦ��0Z�)Mt�d�+x����s�W[M� �B���%Zk�s
��CpZh��)o�,�KE��:�ki)�[��n"�0�U���UT��3��m�hşH����3$��q�]�:��.��4��ڷ&y����q{�-E�)�(��S
ډǢ:�-��需_�b����!T�2�,�D��&������G��\h��(lI����	~讥'��E��YVM�ݠ�	񬁭Fő���f�4��ԍN��/�>#xfE�FP�~���d��e��3�z����Q��wK�
�6����L�.��ቹ�ng~1�e�"�өARm�z�À&Lg���:�؊j����/�
��3�Y�I#k'NߩF���f�L�=��i��L.��z���?��tyq�d�6��ʌa�A���>���Q�/�j���T�Z<RB3î��N7-��������ݠ��H�ۤJ)Ա�'�95���u���shʶ����ՠs�*'`~P��<W�1m�QDf2�D�Q=��V�-�Z��g��G2�tR��./b=�~jr�ɫ�2��I��k'F�Sg�[�Id�to��|	��iB[�a&St���S$>7)
+�*o��Xs�`�|wqϚ�����^�q��å+�p\�5i�����$�ܢ���:\t=l�\�|73��b���6Ę6���ԙ|�s���m��j�#$�U.ر����>Mp���e�G}e�n�7����m����;�8nC��a>�3jZ����<����@�ݶ7���t�#$ R��fmq G�㎲�M�����uZ˖��������!m��@�^���։�O����4H/bվ����
���li'��;�;�є�����`�R�%��Q���e/���pppk ���aK~~�6��E���A�_����Nˆ�@�j��թ�9���E�3����ڥ�¢�����^d�I�9оY,���U�h�drݩ�/�e�9{�.����	�#[a��Ŭ�N���U��HDd��L�t�rY	m��d�S	��FGER��Y���l�jEz|n�'<�͗�5����WJ�ͺTO8������/���Jǅ��S�0��œ��r�|RӰ�:��c}�zfj��HA���曇�2�C��J'n-RbjYu4MR�UD˓_,��ki�Q�>9z�֌�-k�qA[anlP �Ti�	�@�*�T���n�2��t�0x���'#�s���`��DI��3�����}���o� t���v�	�P����g3#�XiB �6>�ݹ��/���sV�9�XAI��h�CX:ܰ�����:[�8�Rw��,�������Oh~��y{jÇ��t�ĸ�vd�a�w1D��t~�p:B���2\T"�K3��E}7�6���t0��mq���}S
�/i w�uy+#�&����������dF[)��./�������h���9���o���s�&1�	�JT�Ќ�%��K`�� ގ���&��?�l�H$J�tC���u�vy�#�*?~�u�E��5�'���;�b:^_�w�����a���7b4}���_9�����>H�{z�BDl2Gp�@��M���3xf;;�܇�����&�-�2����u �6��DL�
`�3H��^�,�/�W�LЈBkn��L����鯲x��l�\:�~m}�	��e�H��D'C�`�Ί�xM�3�-a{%E=r�D�	]��:pK���	���j��Kj4A��G�/�S�?��L��X���rA�5�LҔ��I��5w���&�E�B)�� �+lO��m�"�]ۇ�9Z��Ձ�ܒ��>�9�2����7�aJ�-ƽW��j�˞���qp3���>y��.[���c�\i}f�wd�'���Y��^䔙��qkb�L�@5�#>X��'����['N�,T��8���oI�'�H��߸j��	�֛�)/���ys`ܗ?R~k�X�
�z6��X�~Z)t�jza@��8��D��Ù�e
Ң�9qR�Dii��\�wo�n���b@؟ 6�ʙ�)���@�!����~���f=�"������ #"t�E����E����|�(���
�L��3Ol2�@����\�ɟ��"^��
^�@9�_�����o,�d�o�K�"�/���d�ԑ���KN]�d�؄�H��X�'-�z|	$���S1��~��&%%�P� :���Z^�+fp���7?	� 	����\����uL+.!Q�L��,��h��Eq�hoeE�a+�?�m��'sny7?CA�pE�םSS�):�"	R�/)����܌�[B�ڎ���bg%^�(�X#e�;E<�2ީR�]�~��Z�}���T
�(�O�V�Y)y�P�
_�m���f[i6L�;%�g����Z@ҙTH|!���%�
7�!� �o��
|H V���ԏml�a��%��;M�����$�cDt�=�3��<o^Ð������sVa�!��+@�޽Z:�9=J-%����;#��>8B�ר�|�gٖ���1�&"��`{'���z��MJU(,�п����4Z2��W�����7w'��~�7���{��� �)�nW����#�}{y X�tWZG��1�F�(HK�����w��g��}毱�ܸ̰�)��d�u)b�Z�Ԯ:݉�\/\}J�9e�ꈹ<eQ������5(�_��a�ǆ���4������d�FV���PLVG����TI��� T�����כ)��`��?X�]|4�f띞�5�� ���w��u���S������:��D�>��,���N����<�����GFy9���	 �s��r�c5r�ƿa�8�µ��=Y<4��HL�"܀y���r,\_d$U�_��Q$�A�?����xq�43G|Zf��Q��{zQ���R���W���Y��t����b��q���@m��ݩ����Q	����@�3�d肂���*���	DN��v��p�6ԛ�H(� �V�O�6(����>��A�R���A�c��-�L����u�j�]��E��_�8�S.��f��������5k����*)X�D��Z;����x�(F�Ҩ�J���mkm-���{�p���Osb%�e��s�hd3!���$�u�
������p�kms��V<�ySNdb!��	�x,��cT�3�����aߞŐ�Z�eTPL��8P}����E�2�N��N�Y���9#&�ř�1�������s)���T�@c]Dk�Vh��R|( @�5>�b�T2�n�l���U &�f�iV&Z��*�>d�v���ad��G�W:4Y��f���j6�|�Be�<����ϊx8~W����?wD!i�R؀'H��=m�n)ɊrYi��%�6*��v<��W0k���r^�<����4�v�	�?yq�+�r*V��K0����0�M�˺���n����j�g?�=C��F�������5Y���V�n#���?ǋ�{�
e�۩�>r8/c˭J}w��n�"U��|کg� �&��*�dK(<5�����o��סT�ѹ���h�/^;�u]����Q�X*���2�V�v�l�A��������D������.��X�ڱ��4���x=���:F�Vf�-9�],�y���$�ʬڦ~XoAVk92��(�%B6�h���o�]'�nD�!:&=v\��0�j;�`�]���*e�����,<������Ҭ���zAݔ�qR���T>��:�nfa)�<��\�i�:l��� �9B���|O��ö�T�$�V��� ���T9��G|��f�nH���Q�Sl'�8W��#�r�pL}���%q�(s2;������o�
�:\��x\"��]�9;O�NKqN�F�VP4��()VX�V6�T-�X����ْ�S�Q=���G�^������u@Ӧ���f9yQ�����AZ�ޓA��2����Fe�4P�o���Va����		��]�FD�ʲ5�ro�W}X!�;�i$|�ؘ&ֶ�ܥy�4��'��S�v�+3#�郎��W�����~2���8��FW�acl�V2z��h�w�E�`�+|'��M�����/�a�܈��^7������I�'���a;1��wn	d^7��~W��ie�ѣu�V�s,[x�\�x#�?��.�m��*��WE()��>Y<
.T_�gb�F��q�\�0��J�ό۲���|�rS�(>5b�R^1�SW���5F�ps ��i�3��30T/�pa��dPlμ7�?���M���?�-����:��=<_�����$]Uɋ��:�v�}	�3 фW'�l��.�����sJ��YO��Wm��'^;e�-�9��r\�ܶ�}�W����[W������#��HL���5`��DŲЇ�\�O�2�PO��Z�E���9�"T���\`���}�����tE$tŏ@�!?Y
u��4Bb�
[���<G�4�]=|�>MSF^<LW�z���?�=����
��&
�!��W�O�*N��-{|P`&i���"���Lפj��9x)�b�n��U&�Ĺ�	��#���|Ć0���k�\D�4�*/Qlb�
��-]��S����;	YD8|�F��a�����tS7Ҍ � a����4�u{��v5mE�#�}x Qb�6�N�og�
'f��^�P�wml�6��.`<|ܤR5ɷ[��ʹ��R#�.���@6Rz<���Ǣ�c�����cNk�7��U������y�֎�S��h��p��--��H��A�=G-m�uk�K�X9n]�5�m��ʪ>�~��D>^�3�J޷ �˫��~e��~�}�b.���Ζ�1_I��)��B���c�.��K�	{�L�싘�U�������"<�#|n9VbL����M�ejo���x,x�s��n,�FH`�L��u��B���A���.����
%:��%'H��@���M���d�ٗ=��tj�*{�y`1�	>�t:<P<�l�JЎ�"}���{�8^�xt�a����M��7�
3C:�U���*�D=�Ƭ��*���Գ��(��B��q�����%�VRr���*k�R3 �oth���H������֭�����C�q�9�l���)�;���C�9B��Ȑh5�SG�{8���tњ� �CK+ewS����;b�E�\���A�Gb��Gb��zǭc����\��t[�/Mx�H_WǠ����ޮ7x}��a'�w���zWU'AtS Nhf����l[��ד�l-�U��#����������Jm��0[x>�!UJ�Tx�=�t!�]��HֆP	r���z/��S�,�b]�:D+�Y{��4r9
��֊��	�[3����k��|t��~x��ڟ�<�-_�ۍK��5u�V�8�^;��H�Ŗ��u��
�^�t���>�	3oىd��^(be��54�Ps���tE�@�y��m���T��9)��k�+E��7�\��
�B�:�L�����t�	���+��{M��q�Fw�����B�"�K*	���~ӻg�n{|�Q���Eq�^{ϟ������u]QQ&��������K\���Q=dsws;���L��:U��(0ob*�U�����,\^��z�Y���lt�0qL�?4���+/�-�7����^�4~-�XK~#����F�--����^��H��qga'c{)��D!�$�?�kc]J�])2���S�,Ҝ�aaP�_�n�Y�5�Yߗ�r�ϝ/�|�'h�������˹X ����9���O,F�F	i׉�_ϧw��	����
U�$��F�� �\[l���~vtT�^�3��I�r%mk��R
ʼ�:^i�.%�!�f��!�b;w�Njq@˧˶UT�+�D@=��Ͻ���=��_�!6if��}��hʚs�źKJ�#�j6��B��|&/[|<A㝳�`�oG3����#<N��pm*@�쁄'���
x���:$��Z���8����!�4���{�)c����^!"�;8�Ɲ
������}(��;�_��Ws_,�1����6!O�Muzq��u�J�ip'1�pG(��K@kS�! �؊�=�X����i��EJL���{�De��;-��҅��uY��Y����)a%q=փ�1�J�.���j��w�K��N�]��|�|���y��m	�M�n>��N}����B��U���E����|L
.O�Y%W��,����k����[�(��������QdKq��U^\�M}���)�:�z��	^]ʩ!���Mb-3pE�˴�^A��b��>���v7�w/@�qu�с#��o�6�;{��N�K0�Vb��}c�Q��u��W���f���VdLu�b?M���v������1���^K�-aǍ]��f���Y�y�1݉e���i�L�U���>qd	K���eu�{0?���a�s��M�,C<@y���V�o���Y���f��"N*P2d��$&P�֊�h��q�A�j��KlԿF���"�=��g(�ˏ=;��ߍ�&�<!$bKi"����'.�������h�튍X�<�ԜHi��4� =	L���)����SH°2}���=��ʴ2�6����G�5ѰZ�����M�S�uCxt92O[��\�)7yB�bz����k
��h&�o�lL���4C	0g�d�X���/;m��Z[%���Y����*�T�ƅ{�'�R��.���&��u��R���s��a��h��s0��s?fx� �>�{Ԏ8db����C�Z�(��z"�=[��8��B���*��֪�WOʬN��s��B�3�	���J�8�8����4ژ�˘�R	ܗE�U��(SHԌ���gd�crt��`$�C{�m��T=�tѰ�Q���"�Z,d6�E�Cý�f(e�U�2T$M@�v�w�����M�n�1X�����U����NǠ�vf�<�G�Z�n$>b����ԡ��l�DSa�pCC�P�3cw:���Rc����e�Ϙ<����f-�)�܁?�SmM�ڰ����_�CDYjLS�II��~�Ha��aӉ�@�Y��\�J�tS�i�9����0L���8��y��@-���w�E�1�h��TOX�IS��z3�@�qO����vˠF\;���x�m2F�1����U�qC���k��d�#q��}�`$�=H���<׳�^�䠪�uY�BQA��P��� :�`�S�u*4�.�������x댒�����zߝ_�\VT��}�p������y"���	��������>�`����D5����o���������:Þ��4�ѷ�H	:��a��z�GQRK}k`ݝ��-']���s�)��^�x1nH��w��ùۂa67���+��ŷ6�#jj;��p��o��7��	Φ����t�%̓���nj�ӳP�Z-��@��]y�9N�?}��J�M5�(��	aTH�A�"6#��!�xẌ́�F��$�PYs@�v���w���*R�e����.��W�����Os~@�)E����,�~_�1�L<>��8�,�������J��X���ꪅ���&�Շ���>e���Ea�:bj�È���E������?�N ;���<�t4EP��s����FN=�&x �U(;��.�^Z�D�ѯ���[Z�	B!�*w�Z���7��mMg�%��6%@�yl{�-������S~�^���"�2����3�ٸO�O���N{��27�*���,~ �@F��K����pٔ~��/���B�EK���K�ꙛ�Jt�Ej;�]{
D��bG=��?�"
g��G��Ҭ��}O�P����J�i�����#�����Xr�)vB��s��X6�oI����7j�n�d�O5���f��N��B'�}>^	~�h1j�)7jc���u�މ8ӏ2Y��R�  
b�a�:�.�%V��!�y��xB�E��a��� a��mBllh�X`G�]�㳕I����*[�;,�0z�T�`�dV�:�œ�9�S�|�����}0d>������|��G/jƼ��7ߕ���.�t�nm���O�]��C�Oh�ȡE%/ ������������ͧ�޹ϫ�(��dt��)%9w%�#qu�ؾ���F�??t�����}���/��Lt�
�u�"3m�Pϑ�%��T����q?��[h9�hGS!����2�xl�:r�^c�TUf���}����6��3�	��̫l�=�-b��q�]-n�&X�t� �)�������j�Յ�0�y�sZ�Y0ՏW�糅@S{�ĒW�ko����	�nx\��&�Td^��W���Ρ�g�.6�ˏ�D�H�s����`{��P\ ?k_t�g��J/��J~��˝�m������0�r���X�@�Y�1�j�֜ϺG!��ְo�u�(��3R=C>{>�`�o�|���Z���Uz2%�����^�X�� ���'���+Z=Z`�����tq�0���B���/8BX��qq|��O�~���Bm/�0���Fr�n�3�N�t��"��}�/FRG�AKD����s�3�|@�fzHh�7�W[�]r��w�������}u��}?��֬hЙ������&ȧ3����j5~�Mᵋ0�R� ]��˝��c����(kjR�:C랆�ӡ�9�@k9JRy�o�?�M�6/,u8Z�R�v�����ܞZ>wE@:��H'��S���b*a�'s��:�;Ĵy>pi�$���d�e��Z*�S�:e.�ȷ� �/�0f>(SN�EV8��a��;L���$7��+����P�3�Ƿ;|A�^\���(�<�e�=	�1U�;�G�!�V��]/a�%��N=��/КR�R��}ρ�@3��,�O?����oUm�'�:vkv�[���J��-��^'���%�x_���w�Ƨ)D��#l��r���N�yr��8>\oKc��$~H^սdđ6�����b���3H��ƽ>�:TIC�&:��{5��O��Q8��$���`��������%%$oA~�d<�B,�t�ܶ���=�?�<iK)xC��A��9�S���z�J��j�2��O���G1p�}]�-öʜ�e��j�ֺf[�Z^/��_���
d�(�4�r�PJ7tu9#K������*jmկ�'e�i~�*W�ɠ؉-;�r,:,�,l��$N�Ծ~�^��e?��F�'�`��i*�6����r�'�,���Lif������s���2u(u����1�i Mm�S�θQ墣 m���~f�]�g�뿃 �(ֆ�7�ڕ\~!�g)F��I�T?Z����S�xJ&2jB�h8�Z㬽�d�i���O���D��yS�$�:�]�X��'w���!�e���#��˴�*�'`��7A��53����k[���F��ڰ
��������h���ˢۜ'opv l�B=�c���8z�E����K�Sf/�_b�&��J���߯I��
 ���>7{cs�gIK�h�^Ղ0XFA�Չ�A�q�3/p7y��<j�^p��U%���R�2��RH��K��1&����>��m�	��-*����D�w�y����OZF�I�'�/�|RI��n��33!��f`�c�s�`A{D6�U��p2��Ji��+:s_�oc+����6�� @���h�xIY|ˡ_�41�Ě���8t��׳k�o�,����,4���W�4Vp})���b����P���.Qnr��	CI�r�v{�� ��ބ��f�Q�uB�s�T�[��]�/s0.��D���)����p3��=F�$n���_��K��y7(�]��B��>5���u��gx�Zu_~���H���O�Ɓ�,w��cl;��f�����.��qg�j��(�c���6� ��[ ̧Cc��t���)�%Ά����t�[��[����5�Vah��ݣ�b��޿��_)�����w����xg��9�b�8��R'}z������� y��={�� �M�}�W`&V�B�d3 U�_���$j�����4�~�v���'<'�T-��A��xd҆=$rY���Ch;��4�m˖϶wi ���Ѫ���Bܵ�b�� ��>X��P�Hk�"�1���q�ʍL���X�ϭ�|d
�*@\��[�k��h����VR�4^
�����y_�"����X]J&����8�f�q+w�]��l��%E���e/�%7�����n���͎0��8;&��K����G��թ@���[u������ ���)'*���&��f�fVun=�Њ
�����܏����;�k�]�|��y����3�
�W�$��������+h�Lpw	n�.Np�݂������sqww����0���5��Z�0�������ڻjױ��{ֹ�t�������x���B��ƫ�����}�_�%n�Ų����ۀ����Ҍ���G`Buk�43ݹ&��+�ڷ��ڽB���Α��}�bY���8�$�9_n��$xܭW��i.�����m��,���qH���U����d!.#�ï��]�s�9���Z���5S�H'�!#U��l]wZ����]�$V:IQ�M���z�n)�dG��ȀS�6��Y`j>e8�&�;�Ѿ>^��|(�Z�ݎ,���R��N��i�{�;ᕈ�V�U�l� e�N�i&Ad��\�u����C�?�㰃��k�Vm�Ϋ�9�
����O�~�E����~PYE��F#� {�1����u�����������l�Y�.����i>�Z
��yg����(���4�f|\�3کk]�lJzVH	�z�s���<o��{c�c���;$�a�u�j\Ҩ*U�L���k�md`=��j{�¶���	c`	�A�������{ډz��s9o��Ͱ�yc04EU:��S�*��A�A�z�����~!غ�)����1�䮇fB�"�x�ѽ�}�'1>�-�����v��8=1���Gco�gF��AZ>�EH����='+���q��"���\{}&�c;�",�w�L9����QXe�6v���2E?��b-���_t�$��"s�?�vÞ̹:,ȅR6��C{t����9q����l_��f7ȉ�7U4���=��fۘ����\��»Q0�1�8��Ю���0�J ��������%^ýkʯ� �r�Iu��uW��Ic���wk�s�h[	�4	g�w�^�������8���.��8)��?g�(�<�_@�~�����M3�����)^�z8����AP��s����
��	����Z�pl,���|Bp�2��wWn��+z�݅ug-�A���5Ԭ��%�[�sB_�6��R�8T���jA��OuH�eƀl�8���FD6�	����z1������R/�^����;s�{y�K��4H�c�9����F�6͛q�!�IQ�^�(ڙ+��C��0�����M{�K\@��,uԶ#�. ,0�`���C�4g�y%K��H�=wC��0�Ú����*w׬!ܟ�����AnJg����I}S�����i�o|I_�{gu��QC�0\�����Np�ϛV`Χj��E�ҏ�a�|y3S��u��Y��"s�e'=�;n}&����9�2��[�8NW�ڤ���0SO��݆O��.=|�D���6 5���c%&Ժ'=}إ�U���ҕ�O���V�����C���t/K�:�W�S�N�hVF�!�K�QĥŮ������̾�_3r7��wٝ�q�����u�3S����i�u�)F�)����>�-D���B�,ME���S�sZg4G׃Sv���l��l�x��P������t f�;~ ��bH�6��J*V����0�e�4�f^`�ڠ���}+�y���f���n?�xp�u���1��χ��ǖ�@�kT�َx��ni��%���>1r����s�c��<b>��m�61�Kܠbq+�n�����O�VF���Җ_�Xh,U�2����r[G�Rk:||���.�-gՂ;S�`�ǆ��k��;.a���k�a�t\<�#����ם�*W̻��%V��" /Sk���i�snU�԰ż����2����ёҷ��*����,F-&l�� e xwy�01TD؇�_m�K������،~q-Ҭz�l�p���a����5�Y?T��(�s�Z� ����{��y�&��.�g$XI'1p;ּ�JE��IB��D���Z�|�u���(t�w/G��J*����vGD�^��T��0���p����ji�k�,�09?��5�g��;�)�.=���*��� ]`S�S��]%)~J;��}^�~�(�S	%���G�摤c��Jmw�t��t����G,{>����K�5��;��!R��_�ȶi;+4� �+�Z�NB qg��ּJ�ui+ |ek,GQ�ޝw�����h��n�0g�v�T.w���rs�>
�V'�۹�E�l�� '��Q�
V,N���U��`�EԽe<����L����Ի�!t�Ƽ/Ѳz�0)w���}�CAL�V9F_W1Z+
F)�*��0n���}��yht�&�y��ƪH�������N�#��*փ�C]l��pT���*�hǔ��/?J?��u�������6��E��8��~}���3r;�nu=8���iA���ob��ԑc����q,����C�L�Q��<�"�N���������H����gւ@,��L'Ʋ� �<���)V	M�R�%�/�)A�2�a��ȝ�Pݙ�����y�S�؉>>	]?X����\�l.��=�u�>�0Mw�p���-����dr
�BE_M����s�]�o�Y�[-;�ܥt����ܳ�Э�U���H9�qiY�ڄ]R^V�f۝�%�7!��	0a��%_m�5j<Q�4��+:R{��,]�S}.�U�n�O��Q@?\�@+��F&���6|.�Ƴ����?̝���Z�&�Tյ�#�pO�.�9��e��rQR{�A��'y}פKq16��
DB%D��t��d�XJ�I�ul���J����)�ص�� m������v«��D���<���R��r�/�鶀���*�3v�V����H0��6�՗���ޓ��Y�����oA���f�f���6^��G����kj�}�~�O���!�G�8$r���$�x�^v���^�T�7�XY�E��4Օ�����)�PtAگ�2.�n���y�W�K�%�uy���v{�(�̇R''#*1��[+<��Niu���%K&ZP9~�=�;��s��4B�!�.C��R���.'��-)HSBz�u�e�I���A����g((�K}�Lų�g����E��V��osՁ)͂��!�i��%G�W3\����n��Kع�u�6��k��蛡H.Q�Q�>��\�l���� 8�/�K�/�L�,�)f��,sB��YyZ����@(��R�x�R}}��LM������HH�
���UnΫN�ap�ӿPb�tK�O�&_?��S0�n*��8�?X�FR=��ٳ��ھ��!ޠ���}�&/Y��T�y���������=�?(3/�G�=/.4w�? ����/��6�~ù?|��V���p��[m[��Ȣ��j��EqX�c7��Y	6�W���J<J�SZ�Q�(��1��!��r�k�c�w���S�䞉 '��;�Z��3D[�Kъj�n�JS�����#�3k
Bs�|t�)�r��s]=��S��1��$��#�d7������i��3V��n��pj2BWmP�s� 5$T�nXV����;�r�������iE����o*g�	���1�2��&���x�?B#z蒭)�^`e/�5d1�*�FGsJr�w�]�m�'�����&��8A9ˀ��]ES����Y5�tU���=:	�c��(�ؿ�F�ڪ�"��i�����J��d�H斔v����Tg�Zc��[��� Ϥ�VIFrz������"�]���R�ѥ"D��>��H���E�9 ��d����k7ڕ���t�^����'����PB�@������ؔ�;`g�,�8�ƓC\���|t��UQf�E�ː�f��֘{Y*q�*t�<����M���ѭrJ��i�R6��Ps䃉��r�t����w,\����oӰU��a�����oA�)�{�%�?�>P;>{,�O��3,�6���,/br�f�GNd�Ќ�+�$����RGp�D*�;�Q��O�1�E�j���a�Ʀk��'6ս��w)�������=a����êW|�n�;B~�`�,B"|ҭ�K��m�)V��O�p��
��r4~}M͐�7�Y@���E��zjQ/^����;T����9�oo?N�U���&ew`�HG���1A.Q��I��cc�
J�t�ɪ lP-�YvE=�J��k賐�"ҵL�^�,WMUHQJ�����}��!��q
7t�����0����V�����o�?��:<�f�"�+���#}b���H1г�� ��W7�f}��$CcW���>N����< �p��}(��9���ɚ�S�K�/'�!���8�rVV�ྒྷ#�+#d��O��<�-����K&����j�wm�ۆ|��F�=�>�]�����C��O�'}}}5��4���b0D`��۵�:$(Z�6c� �j�p�L���������3�����������2��q��3j�X�Q�����&jkC�����Y�� ���C
i��U;��v��1���֤�H�<n٘�T�����a��1($$?7���J�6''g�+:��p9D��H����ϟ����w8L������YeA��:.�I"Z�&Ώ���`n՞�������a���-�Й0p�V{
�K|S�=�k�CC���5!�fN�bn�S�GC��pxoow����7������&H_�?��e������Ē����ԛ����o~<�.Vi���ة��C:��,�|NKK�ҥ�������}Ɵ�"\"� �֌����2�[�<�ި�րC����2V�����$��j9O#�Ń��C�]\������E�Ύm�q�O^X�ӊ�t45X�ZQ�qg��v;�~X�9H�g�ebd��z� j��)T�% �u9��E�^m�����=���������
W �q�{�E����� �ѱ0������-P��뮋(=h��y��tk�s�����3{TX��rI>0��z���(�8�eL)�	8Q�ׯ�{�_NJV��b�WW�Ηk!-,,R���t=�w��t�L�?���l4X$����^4�t���˶y�:��Sn�uѩ+ңT_e��6�����K��P|�J�QgK�����$qt�N��3��8�ڔj��Z���4[�ɼ�	쬭���FEC~����8 �����Qы.�twvv�q5��'��~Q��)���.�\��i7�	ä6��K�h�z�of:ǹN�����?[��&�An�6@ϲ��p��K{X|�{�$FHDV���6`�3Ĩ9h�H�l��`n�*,��̾�<��@+Ms�;�e0����\��Z����i�3g��?���� ���(���*wo,ZM8��c\��P����Po3n�r��A�3ێu�xa�7}���{�ީ�B���ۆ�S�Э�aX�W�پ�
�a���p{�s�>��^i�	�Bں��~O�?��&%w2�g��N۸q��̂��vx-�ج���L_��o3���~��Mu�����c�V��&@+��Zct�i�3<�{{rX�8�z����TSv���\�9���i ���{���^�ކ��Q�#��j�[�8���yj����~q��&�#�qV��W���F��L�s쵘cGj[����?��'�߼Ħe/ʌG-��d�O������|ן2����Ki-���桼�-��a�^���G���553�7��Q�yB��H�����L�l֚X⨶�X|^�P�1n�����H7�/K�eU�[5��(Uc���xs���wB}yM<�em���Et�}�AAy���-�`=�쎻)��Ά,�-NL�{�zӨ�/՝�wZ�����g�!��c"@���gv[�e�m�="F������B<T���eI�z���̐�n��Pe�31T{`~~F��p���y�t��
����`��
*Pawӂ[�{�J�ɻ9vj2�SΜ\-y48�[�zF�ӱ{��_����Xv�/�v�E�����,JmX�&w���e���xBv��受�+�~����,$'����нJ��B��A����l�����erώ���T�e�3_L� eߙ��._h4�'=��MP�4)$���]��S~2����֍7O�k����J�xIX��P�D]����������>�!���yF^�����@����Ǜ����';VB� /�@��Piv�GN��>�ݮ8䘛_7&?O0�cO�H�o�א�N��:I5�%{�sVEy�����H`���ZxS@�R��R[���p�֨aT���&��5Ƶ��@�:M���5�9�Jj�]IBn��:OC��h��71@��-8��)u�Z��G,S�M�Z��W���G]��[��x���S����[�]�O����Z��l�3��5��7띖Z*@�Z��Z_p���As+:h�쯗�yTX�?m�=�4E�,�����ѿJR �\����*�UM��I6g~ږ5��A�/��^Mm���2VA�R�!��q�z��}�kzF>��G2V�[��5�t��=���~�E��I:;V� �%+-ߺ��u����cp�s��۽\�c4��$��9wф��O���F�gY�oxz�7�[DZI�B\�P �.�;�}�
�����*�k�nwvX�1�,G��ɤy˙n�w���Ȉ�V�	�>�� ҽ�}��w��J�"TU���:�8\B8�j�rX�?�\|��p��w;""��X�T9�5>`j3�m.=���C�˻����VT�XH�+)O�.iG?]v�K����Yi6 �n�EfW��~�lC!�ɢ_+�S��R�lq |����[Cԯ�=�u{n�gN��s^�7�d��f�Z!a����R�^��^�������������Zҵ������k*�ŌIAGx^���P`'���p�+?Tv~uU7pWWf���:S�Bغ������tX�2�=���t��&<�������,��|[��4��%ԙ8�k�����׸;��p��-�uݝT#�﬍DIJU "@9xs�cRf� ��B��9Џ���(�ꆿ
a�w�VV{��i�1��i�<�ibg��f�go}F9���1*2������x�c����r5	�y�y�x3e���3'�t��X��v��~h�@<�����!�|W�IZ)s��@i�KOޚD��������f?�*Tp�z����<�8�=��\k<��.,��L�Ǆ��p����R3�;ι¼�'�!>./��,[���u�a���tȚߺ�oS��s��M��8Pc���g ���|���ZYCfS����(��"E5e�mCȈ�}%��E�}��� JU(�䔱�&��P���d�� �*e�h����Gu�u�t�+kl�E�L�y��!���9!���`�/e�̡��y�U��X��l��_�M�4�v?QmDt���2c�Ldsӧ	�W�j����"��b F�#4�_|n'%R�Z��	�M�Oh`٣���\��=2��t�"���n:o���iF��1�����$/�=���;��@\n)pu7�PT�$�y� �������^>(1�ĔCP{��z��HI�u��{�G�Ę�����]��������1�X;���MU)�ZZ�B)���%YJk�Gb�N��	y�����<��]�(E-ɒ�R^� ����x��)N_\�J�Ɓ^�ݴbi�Y��k��n2���l6�[�R�_x|_C�=�ŉ3k�eKSYE=�m��G� �������E�ƚ٣��?�'d
L0����m"���Æ�/�E�9)�:B�z�����b���P���9���^������)P�	� �G��r8�[Я9уy��U��6c��QM��� Ր��p˻.G��{-�x�>-6TG��O���Fo�đܺX��[<[�S��$�#��z�ܚ5=�\Ҁt����&Zd=آm��rK���G*��}�c���\��:�Wf�p�/}��p˼ص|��>�@��ts6��Ix	o0��i�Z���'��^���z~ �͡������0{��s:i����~w_�-�a8���@�yJr�}�H���{�H�a)�Hw:#J��/�K��Q�b�~8��_�.�5�i�c&*H7wn��?��%�kS������ל�2��e:Q�.q��� ��U{��p�[��߳�}��G��?��~U�(��+p�̲�<r���IK����4R���\�[
�I��)n�p�Ѹ�S<��Ԍ���W���8���0�iz�@�����%X�
�xޣ���-jЙA7�ɼC������h��D����tЭ+�6�Ϭ*42�ݒX�F�~��>gˎO����P&�]w{�`�.?��,���Kk�b�_^:VZq����z�&�«=:,6��?�X�7ɂ�(�3y�Ģ�gl]���pFۈ�<��1'��N�?{x!t��Ҩ�Ъ�V��:��2�MWq���-��gs�<a$%��"�����(�6��*���=��,��1>6����XsB�ޖ7>��N*�������M�z`�p���Ǒ<Gm�OA��Va�&6ӻ<�'�~{.³���f�[����el�&t.�I��F��5��<�r�,�n�c�|K��>X�/�����/�	ł����kh Xn���]Cг��C*L���Pl���a5���T!� 7j#ǟ��J���ϾX�g�%��<J���*c��o�����B��[U�!~ޭ�-�,���P��!P������`~�^�w���/��	Y�q�Y)�ҚR�����9�Zz[9�T�#��_��I��3N���@ʧisE�F�ñ� ����5o��X���8c�\�\`����~�D���Sx�����חxn7��ڧ��t�֜l��SG�_��ԛ�j{\^:�����9�{�t}l�[/j*���~h;�I�0�{o�6r9A��뀭�g��5u�=�Pt�gШ�ڙ|���R�OV�~\	oV�]7t;a[FK�qz��
�	>%�5EE7���3O�;r�>Z�X�N�Z,��V��߄�Em��S�R6���*���N����f�f��u��n��� a��m�ʋr{���-�ݯ�7�A�EA�����������!-��Y݃�a��[V\�B��&����mE������:�&t����u~,���A3�" ��j��Or��{�3�-�JB��w�u�<&��:b��ýo�߉*\s�ER}�پlq	�7�B�[͔xau}�&�}�y�y2����~�a%ê#��a���y5�����&6K�"�S��a��fW�J_D�ϡ�ӗ�`�e���0��uø���L0��l����g7Y�R<�hAwy�[�{����7�	Wm{\���m��[;��k�^��$���"�u���Q)�<Ϝ�����P�aO������y���T9�YB��o�'�	e�l~OW�.�G����5Y_��`���P�u���շ7o=�ʰ؃����?D�/{E�T�WҜ�9�Z�锫���z�'#t^y����r���� �Vg*��Ap58F֓�]��Q׻i���P5�;SmhJҾ�\�<��g	�Ӧid�7����dK�\��Pr�ԗ	_4����髋��ݽ�?��9�ʱ&�o�󗝊G�+�%Ǜ&�[]��w�Ni��7E����F��A~�ْK���P x4���}���x��W2c�.���3���������˛^�U
��BF&�,b���2�|�rf.���/�)�@�UiX��nʔ�.��?������7��Z���GKk׋�iֺf&[}�����;��?gX���D�N�[:X6� I�xF�������eK����ۀP/#5;JqW��D�5
�����E��}� [1.��ߪ�G���_Gؙ�t����b&g��n~84K�m�89.��5/2�1͇��L��3�G��G�jqV�\��]�tvcA��0��^h�F��qF;�}������a2(��$�%�������%o��|�p�R�O��țoFq��|�f�({���E���Ƒ��a��*n�L���;�yہ ��]��R(��3.����s��"�2����YB@�8j"�?%�y��h��l��t?�Y��>b�N���7�s ~�Ei@��`��R��U��V�)��j4���x�R,�#[6f��)E!k�(�0���.��W����kF�Z��1���9������>�IZ���^߰ )�&���Aݙ]�--�2`��>kM�BMf��$.���N�>��a?�8�	c���~Q|��h�8PS��0N�#~�f����Dm.j����h�+�7����i��[�ܭB`�F�|P�c�7�x��Ln�Ӂy��@��
Y��_�N��k���%~� �My��j��%�j �^?aO�������~���|����iZ.��白���V� ���Z���{2n���Q�{|�xMz��~E��'�c�̀D�ѯ��ޛ�r�A�k��74v������h.=a�g�`��������7��~�{�`��I����(��E�>�+b`�%��4�do��������޶漱�am9����ꇸ�d���ms��Ru���m���[��8�r_d|%\��!��%�HY�)��5ӈ�������@�:��']�O%�����N���u�yi~%�؉>Ƞ��5�u�yj��p�bI���U�8ש%����������'G�8��N�2�[���y}t�K������q�w�OE�>.�h�F��*��i�)O�L���n9I����xi�i��F~먵�R��^7d-��u������jtf�3.�!��&���M���⅙Y�s������W-W�ӨX���(������O1*��l��1�V��`��fG�fNcNO��#я��}�{������K��4y��r�����~�6�i������0�v���f��\|�� -gQ�2;b:��,�JY�V����
a�In�mȒ:*EJ:YD5β�|�\T*��d�V�-��o��x����ǲP�ܡs�U�9V��h<��xЯ6^D:aP�p��U�����0�{�X����+���7pu�*c�6���2���٬m�u����	��LyM��Φ��&d$���փi��R��o�g��j%�,S��P寶y���պ��]�
53]&�N��: iLx�ڔ�Ζ�o�;�$G��F��e�ǰc�Û�V��S�0Τ;��Z�a&Anj�KYV��|X����i;�_w����>�b\�+Vki�ב�K�=�q��>>v�mȬߐ�Q�MM���f�s�ID�^�~�H�/�l7ڷ[�k@=�Ǭ�?���ɪWܿ�U�����K����"��k��N��b5H"��/W��v�}�[�9K,� �INA�y�d���k���ʊFL��#�тg�G�O�Pbm��Z�\][�_!�_���fZ��P�=R���Nm���/�D����(ɡT���.�_����ŗ�y�v�jI/
?���1ٕ�p����n���z,}���3�&�-��f^8���l�#������(� ���G��S��kZA0�z��"��}�$�:ܹ�'*��R��=��E=6�5H�˝`�����u K*�1n��U��#rI����s��sO�3�?Y2[��=�K�#6ĴNQ�<���#��1:r��k@Ç�Z��N�Q�����w��Ύ�a�[�E�nҳ"����u����?�]����,�i�偑:+-GNG�AF�ߍ�/�� ��ѷ�xTf qn��m wb�e�MC�}X�R ��,3/'rQgqm��")\�CPiyfw����e>:�bo���.�m�q�0�i4P��Q�D˱���(�}��0
��S�Ǚ��>VV�ƪ{T�'v̶�m/��_3��>�IEIG�����x��4Z���(�@�4�59�Y��)��r#��n퇜��M�����8m�|;">�B�tI�*h�'��N$9��#3=2�
Uv=�s�y����0Qf<�1��p!V2}�#�F��8�p!���Ud��r��^�vG�8����H������V��r�Yeb�� rw��Qs�1���F�����%����5��k.��o��|��b��K5�ꏒ��ӟ�g�V�Ȝ�{ŦL>��_<����7��7�F��H?��'�z�F�ok���PFvy�)�����,%�ۮX� ���y3ЛH,�ܘi���6��n}P�[�L�2b�����L��B����*n��?�?=X�\��n*q^q���e'o'�PԷ ��@7*�Y C`e�8Y,M�b1y�Tg�|bS�H�oŋig�B<^8Y�Q�^�J���j�g�����ݜ�j�R�Y��Q�a�K�f;+�z�y���jg�����,G�U��W������@��N��Zz�/��Z�TK�(&�k��-���cO��^�e�>S^�o��A�ɹh�f��<07�}?��r������䇚�0	9K�Mv�!���%�Z�`e�����EDE�-��x��$��$���)�7W�nD����#���&�Db�nz�}/z���\��\����ƍ��r��erd�=�kˈb-�Ž����^����3%���AE�f`����6	��Љ����A�mRY��I� ���e=J%Q����~�wv�P�5\� �Ap��tJ;���I!{trI@��Ek��Qu��;��_�Mv���v��T$��͊�B@q0��l�@���5٠��Nro�ͷq�z��q�غ��X�>��QK��Wf�i�JDb���1�K?�U �<[SϹi[׈�fǋvrR����/?��������#5j�fr�r�בD)Q���,d��`���'�����+a���?��ӟ�{�:	�VP.:z-W�g'��U
M�$G64����vٹ�bMj���B�u���%Ύ��vH�vP*��ԁI��rP�iл�p<J����b�,C#�s�"�م�9r��Q��B*|�:�h�a�կ�j�1U��iqV¸��[0��4�/��*@/�'�+���C���~�J���Q}�v��b��W&i�F�ݰ{� �l9#���@V]S[+r�"RcuGhl��#��\���ʯ�&Cv:3�� ����k?��0=>_o(5�����@�CV�E6��a�l7��S�������?!G��i��J�]J�����դ8.�/���-$_�g!���i#!r@���N�$�FM�Kr����������fZ���[߱7�G	�V�5��F�Iޔ�N!}�)'�n��ǝk� ��V�0��*D�Ux=X6�:m\���[�CGl��vo�}vb1�|�E�.Gϩ���+e�{E.1�a�
����|*�y\h�����FQ���T����Q!�9#�?VS }c��F�z ��NԆ���|t�����7P����87Q�W����i�zO�I4���|�n1D9�y�e��|�,��;$%����cn�:N�@Ԩ���q:ǧ>�Ν�ͩj|��:BT_+��
��57�i�,g:>�f�Cv�x�{F��k=_�y(G�O���� ��ҥ``�Lc��g���aF��C�;v��N�<�Yl�b��\]���Z�;�֑�R�j��=U�C	[e�U�ٗr�߿���	�Sw~(�r�Ng��)W|�$zf��]R��S;�s$������F���w�Lm5�P�rp�]��g��(�R���,��$'���|D�!y�g�	��(����j�Ϗ�(���Mv�!���#�\���m�P���q��-��'޻Ӛ=�N+����V��@Y�M���;��ʴY}[�XrS)t����Z�5���ݫp�l�<��Iկ�<�&G�㼼����
�fK��	$�-�
|��o������2�xFط4C�J_��&{�����M�N�T���V'/�J�`���k�B��	F�ҸEslSѯV,-�c@�D��Pl��|V5��Q7�94h��#K�	Zo��Fw�g�G�� \�<�Exp��mI����0#��A�<����	7����i22���owՙ_�7+��_^#W�L�(M���u�c��r=���5D�"���ٝ@�F@��������|���k�A��'�[Z�'�I�Nr�P�{.4D�j �K�2�C�����'��(�T�\%&��J�g9]�~��jv;u��8сv��F��V[MW�;�f�R�M1T3�6R���r9��8[���=�#�4���!��O:�A9Cd��W�1��A~��Ģ�>nϑE��瀍�K~�P�
���ު����=!���/�Y�?6B����efaWC���]`�wK>�E���ռ*9�]�\(��|��Ւ%,��S�}H���Iw��-���%O7+�K�[A�2��vAT���sS�AqL]e���KΣ &�nm�K��)*D9����	3��v୓���:�������zO=C�e{̿��/#�6��h���)ُ�=�9�n��Њ?F)~�,�I)�=*|��f�v�����M��BE=J��4�����̵I���6A�����R�0���uH�4�~V�z�c�6
�_U"[~D��~
���O�-�2�:���&i.kS�|�B�
�0J&(��@)KxD�T/-6|*$��,~�+��MC����³'��Z�[���Š/�Ք -�F�5�r���g�Y�����J�,��-ݶB�G��DV ������֨�4�Yf��I-����Jl�F�a%�WQA�R��3�S�:�[�.ob�N����eSހ˜��=v��3��V��˳��lY� S��4 �0������x:�r~&vF�/[�������t#֍�
��j�]x��9O*#�
Uπ\o&W��������2�<�3Æ�9����i˶�
�	����j�v�dn��K�F�W���:�V��D��e��#G����X����;sy�n�#��E{~�T-����K��FmdIi�Ə�Qш���>+��8���6��UL�AiHV�q(�2�j�<���J1��ó.�D��׃q�t��k����7�<�l�&��n�̎"9l�Vq\�lRHWZ�}�M�"t�/�$����C��V!�r>LG]i�	�Tǰ��=rF�r���l�={�u1��g����3N�'��,��#��N��%����u�E�(�%��*���-�ôL+�[x=�������np��.�6������=�U��r����z���id/�8��s�lY� ��8k/^�%�#6����f3��$��LdL�k M�06K��s�]
�1�|[.KQ�9����s�IG8��7�s��$���$�AX�9�K�Y���@�=#����ν� ����m'������<�w�f�3�>d���a��E��>��U
zc{�o��̱����v��%n9X�٧piGG~��G(�:���L���п0��ċ�3�hX��(ҳGh��D5xj�'��<�C%��V]���A�������둰!<|�n� '�
���"��&���W5����!�i��_�Bт�M��� �hw�o�J������.�E˂
�HQ�'��ȫ^_���Ul��F�?>5"ok�.�E=n_B?-YU�E2U��iwE�ph_�Ȇ�M%4�Tg	���1�0M>@�Z�D}v�F�O���#�J�v6��E�'t?�
|Z6W�[ME�5�(�va%�÷��%��{�:"�#��o7b�V����#$���[�����A:��Z�ɉ�cT�� 
c���aG���K4RJf�8L�e����r���+eI�eʽ ���N���A�����f�����m��t۩t�γ�R��!���L%\yD�V ��*������/xN4��NØ�R��nm��@��2��!m��>R���EC��`R�㻩!��+�����j��k�_o?���-���4�J,�t�o�l�`��H�p�/	j��CD�y��ίԔ���l�ߘZ]�P�}S��F ������J���ܴ�`RP��v�J\����|-��?Q
�A�él�>��6��T�[�z|�-������j�k�>I��/K�o��IA@7�|��p�m�r9P��f㆟�:M㞺p�PU�l��*���e<�����V���D���Ff��.'�MM�}�����i�q�<���4��,>Cz1����YE�\�_U:���'U�q9"f�G	�1r`H�V~7-�N��2�g�"��;k�/����V��uX}�Lk��Rw��Mr�obЋ<���jZA�s<���_E�g�2�=d��8���D�Rs;���/)�0���%����A2�v0�N��� N|�%rs]\���Fs�v��A�.&o�N��ŦR.����qΕ��T�V��u�(�ш�Rl�Y�f\�v�Sq!M�3v8l̈<ig���Tg!�_�$���������
�-]�L(�GP���F��KC���I&-��ɭ�@O�m]�,�P޾!��=I�T�޺��v�����
 ����[��̮u����H��{ڟ�`�PǇ�˝��Ҳ�\y�:����*��v�z����������l�ֹ�zW�wƘ�I
��p;8���I�OP�Ty��XB|4�nǳ��^#t!�t�	O�LW��1�¾��L�Fz���V�ÆHPl��@D9J�.M�aκ�/�GZfÑXN_C�`p�l�gn���	������yU���Ǒ	�X~�	#'�EabOl�3�۾���k�j��e}�hH��阗Op��i�>�*�R��B�2��vdU1��	yPO���4�M��O���W�(�Xh!v+�D��M�B�l�^w��+��Ο���-c��K��T�d�i�7Ҁiu謂B����3�5LFq7e��xr��.�1��Re|��YnnEX�8�zjj2�%�!>�%�^��p�!Ŋ$�Xa�%'���Ȼ C���9{.��+�!�6�ۺD�ˇVh�w��j���ޟ���.����x0���N7z���o��(��k�������w	xp�";�!$ƖE�o��7�Z��e�J��U�wC۰�2��6���Y����.Y-jU`���K��WQ�3<�l1$"ׄ���P�ߢ�����;Ap6_sĵ;����]k
�(��;�>r$��������YC�bM)���B�)k����`�4*�f^/S�U�J+Ą��Չuޒ��E�x�����2�ք���m0�jy���O*J�O���$0���Xޛ�Q�إ��k�9�:�Vp����
G���d�H�������D�i�)��Rn�t�Y($�7�����8��a�4�Y^jg@��_K����J9��[GvS��]J�g��[&�Zq��~;��Y���o������h���-�B�t������x�z_k+����?�/Ii���#}����F@�]�N~�Ss,}���Z��E�p,.��!M�^.���p�Ő��gdf"�]�� E�4<���?ԝ��9�.���vh�?������99K�8�b�H;>1'��k�,ʗ
z    IEND�B`�PK   DU�X$��  1&     jsons/user_defined.json�Y]o�6�+�����u�ZkS��CP�"�u$O��uE��(�+�L�ފ=5O�$�sI�s.y�e�|^��q�v�;��tv|1���uQ����	�W֭�]����e��J�ucY�	9�Ϯ���n�������aG�[؛�qa��9Q�VB�4�2�u0���d���[U�+��]0���s����[���ҭ��X5��ϋ��:%� 
k�r��" pf,�Xh&��WdU��3i��@Kt7M�NB�SG�r7�N�w/*?�����|����������y5~�e\�w��z�ԟ��ү��	�q������Sw�	���f�۲����*gv�ԅg��պ��_��
Fl���� �%#C�~Zf�U��o���F,.����4>���~���#$ 1�H�� ��Tć1|��?}�k���D�¯���e*>��J~�<H c&3� ��2�T�p��h��4z�d�"j(�
���J���W�a��_�d��aGBQ�@����mdQM�TQ��QDe��u��·��F���$L�6N�v,�����\�f��
:��?Uuӗ�	ࡰ�%:��P��T�-.É���>$�h��P���I"<� Yk(�DC9ҋh�J㡘�E��(j�Cr�� �I9���p�&11��PNUSsz	%�T"19�WPY�����s�Vtr�\\�	b�N���y� &����Kd1A'WNrIա���g���M�}��F|*j�����j����7]ǭ�Y�ѕW�����7<n@ܜ��]D��Y� �D�2���D0a�8��`���T�`��Rc� �f۾��o�V � ̔<�	%�f�c���118��߅�b±R8���NÛ�0:���g� ����g����3z{x�
����l��W��F��N��ǉѿ�,�Ї��hO�W��FHC:��]|}v�&�$�x��9\`��H�1�L Č�*WI�a/���y��h1���-��v��MumuEw���vν?	�*4�8��P�$ $�Â�L����Cenq"$(�g��и�ֽ�������'�x�<�p3�Y�ڝ�5}�q����1n@@�&�Y�У����i��x¤��9[�z]��W��Y^-fg��8�I~�e��d�!���Q�ݪ�?>�e���Ruj��6[��V�^�S�{�N��ź0K��V�?۞���n�!:]��Κ�v�޽��J�vc|��=�#E�b#s����
�9� 9F2c%ؚ̉�	��;��D}�w��c���>��]R&}1�ۥR�"Cu� �r�)��T�T�,�8'����E~�(��(�L.r{�.��m]n���nBYvW}���'��aAv�q5#S�5��V��ٲ�>��j�l��t������oO��ʖ��>�R��b�/��t�~-/���~!�AB8P�}x_Wmi}��������9�|���ѤЙP�j��;�9*��fQ���ă@�U�%_��ܧX0GzƆs� .�9���|v;�����W�\�o��y��5m�T�#I/V����eT�Jf��9MM��5(S(�VD��]DOR5�Uq�����f���;�!2�d�$l��߮b|r�&)���&��	�B�r��ҾI��K�HG>��z4<>��C��ȉm�_;J�B�� �4"�L�~�?� J�����B���Y[~��N�?M (��i��:��)�(�3����������߫����?PK   DU�Xx�*�  �             ��    cirkitFile.jsonPK   DU�XK���(  �(  /           ���  images/1042b8f9-2e87-4dd7-a644-1e53cbd80f37.pngPK   DU�X�;�i �N /           ��8  images/10c49116-c115-49dc-9efe-e8b38f603c33.pngPK   DU�X����7  �  /           ���U images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK   DU�Xx��{  v  /           ��Eg images/378c5108-814f-4376-af43-2b942ce8b9a0.pngPK   DU�XH�:9�\ u� /           ��{ images/5bcf48fd-3e7c-4271-817e-97f3eb0e00be.pngPK   DU�Xǐ]zd� K� /           ��� images/700e9707-92a2-49ec-8e41-72cbd6a28b0b.pngPK   DU�X�&�}[  y`  /           ���_ images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK   DU�X(	��I�  &�  /           ���� images/b4edf89d-5842-4488-bd77-04cd2da60bcf.pngPK   DU�X@��)  /           ��X images/f58b3b66-0d3a-49e0-a328-e802f4e45778.pngPK   DU�X��MY��  �  /           ���n images/f7330a66-6727-4ddb-8762-657115be29f9.pngPK   DU�X$��  1&             ���5 jsons/user_defined.jsonPK      $  �<   